// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.10.0.111.2
// Netlist written on Wed Dec 09 16:53:08 2020
//
// Verilog Description of module cpu2system
//

module cpu2system (clk, reset, akku_o);   // c:/users/70735/desktop/cpu_l/cpu2system.vhd(7[8:18])
    input clk;   // c:/users/70735/desktop/cpu_l/cpu2system.vhd(8[13:16])
    input reset;   // c:/users/70735/desktop/cpu_l/cpu2system.vhd(9[13:18])
    output [8:0]akku_o;   // c:/users/70735/desktop/cpu_l/cpu2system.vhd(10[13:19])
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/70735/desktop/cpu_l/cpu2system.vhd(8[13:16])
    wire we_N_63 /* synthesis is_clock=1, SET_AS_NETWORK=\CPU/we_N_63 */ ;   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(13[13:15])
    
    wire GND_net, reset_c, akku_o_c_8, akku_o_c_7, akku_o_c_6, akku_o_c_5, 
        akku_o_c_4, akku_o_c_3, akku_o_c_2, akku_o_c_1, akku_o_c_0;
    wire [7:0]data;   // c:/users/70735/desktop/cpu_l/cpu2system.vhd(37[13:17])
    wire [15:0]adrram;   // c:/users/70735/desktop/cpu_l/cpu2system.vhd(38[13:19])
    wire [5:0]pc_5__N_30;
    
    wire oe_N_57, n2247, VCC_net;
    
    VHI i2417 (.Z(VCC_net));
    IB reset_pad (.I(reset), .O(reset_c));   // c:/users/70735/desktop/cpu_l/cpu2system.vhd(9[13:18])
    IB clk_pad (.I(clk), .O(clk_c));   // c:/users/70735/desktop/cpu_l/cpu2system.vhd(8[13:16])
    OB akku_o_pad_0 (.I(akku_o_c_0), .O(akku_o[0]));   // c:/users/70735/desktop/cpu_l/cpu2system.vhd(10[13:19])
    OB akku_o_pad_1 (.I(akku_o_c_1), .O(akku_o[1]));   // c:/users/70735/desktop/cpu_l/cpu2system.vhd(10[13:19])
    OB akku_o_pad_2 (.I(akku_o_c_2), .O(akku_o[2]));   // c:/users/70735/desktop/cpu_l/cpu2system.vhd(10[13:19])
    OB akku_o_pad_3 (.I(akku_o_c_3), .O(akku_o[3]));   // c:/users/70735/desktop/cpu_l/cpu2system.vhd(10[13:19])
    OB akku_o_pad_4 (.I(akku_o_c_4), .O(akku_o[4]));   // c:/users/70735/desktop/cpu_l/cpu2system.vhd(10[13:19])
    OB akku_o_pad_5 (.I(akku_o_c_5), .O(akku_o[5]));   // c:/users/70735/desktop/cpu_l/cpu2system.vhd(10[13:19])
    OB akku_o_pad_6 (.I(akku_o_c_6), .O(akku_o[6]));   // c:/users/70735/desktop/cpu_l/cpu2system.vhd(10[13:19])
    OB akku_o_pad_7 (.I(akku_o_c_7), .O(akku_o[7]));   // c:/users/70735/desktop/cpu_l/cpu2system.vhd(10[13:19])
    OB akku_o_pad_8 (.I(akku_o_c_8), .O(akku_o[8]));   // c:/users/70735/desktop/cpu_l/cpu2system.vhd(10[13:19])
    CPU8BIT2 CPU (.\adrram[0] (adrram[0]), .clk_c(clk_c), .akku_o_c_0(akku_o_c_0), 
            .pc_5__N_30({Open_0, Open_1, Open_2, Open_3, Open_4, pc_5__N_30[0]}), 
            .data({data}), .akku_o_c_8(akku_o_c_8), .akku_o_c_7(akku_o_c_7), 
            .akku_o_c_6(akku_o_c_6), .akku_o_c_5(akku_o_c_5), .akku_o_c_4(akku_o_c_4), 
            .akku_o_c_3(akku_o_c_3), .akku_o_c_2(akku_o_c_2), .akku_o_c_1(akku_o_c_1), 
            .\adrram[5] (adrram[5]), .\adrram[4] (adrram[4]), .\adrram[3] (adrram[3]), 
            .\adrram[2] (adrram[2]), .\adrram[1] (adrram[1]), .reset_c(reset_c), 
            .we_N_63(we_N_63), .n2247(n2247), .oe_N_57(oe_N_57), .GND_net(GND_net));   // c:/users/70735/desktop/cpu_l/cpu2system.vhd(43[10:18])
    VLO i1 (.Z(GND_net));
    TSALL TSALL_INST (.TSALL(GND_net));
    GSR GSR_INST (.GSR(reset_c));
    sram64kx8 RAM (.we_N_63(we_N_63), .data({data}), .\adrram[5] (adrram[5]), 
            .\adrram[3] (adrram[3]), .\adrram[2] (adrram[2]), .\adrram[0] (adrram[0]), 
            .akku_o_c_0(akku_o_c_0), .oe_N_57(oe_N_57), .n2247(n2247), 
            .akku_o_c_2(akku_o_c_2), .akku_o_c_7(akku_o_c_7), .\adrram[1] (adrram[1]), 
            .akku_o_c_6(akku_o_c_6), .\adrram[4] (adrram[4]), .\pc_5__N_30[0] (pc_5__N_30[0]), 
            .akku_o_c_1(akku_o_c_1), .akku_o_c_5(akku_o_c_5), .akku_o_c_4(akku_o_c_4), 
            .akku_o_c_3(akku_o_c_3));   // c:/users/70735/desktop/cpu_l/cpu2system.vhd(44[10:19])
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    
endmodule
//
// Verilog Description of module CPU8BIT2
//

module CPU8BIT2 (\adrram[0] , clk_c, akku_o_c_0, pc_5__N_30, data, 
            akku_o_c_8, akku_o_c_7, akku_o_c_6, akku_o_c_5, akku_o_c_4, 
            akku_o_c_3, akku_o_c_2, akku_o_c_1, \adrram[5] , \adrram[4] , 
            \adrram[3] , \adrram[2] , \adrram[1] , reset_c, we_N_63, 
            n2247, oe_N_57, GND_net);
    output \adrram[0] ;
    input clk_c;
    output akku_o_c_0;
    input [5:0]pc_5__N_30;
    input [7:0]data;
    output akku_o_c_8;
    output akku_o_c_7;
    output akku_o_c_6;
    output akku_o_c_5;
    output akku_o_c_4;
    output akku_o_c_3;
    output akku_o_c_2;
    output akku_o_c_1;
    output \adrram[5] ;
    output \adrram[4] ;
    output \adrram[3] ;
    output \adrram[2] ;
    output \adrram[1] ;
    input reset_c;
    output we_N_63;
    output n2247;
    output oe_N_57;
    input GND_net;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/70735/desktop/cpu_l/cpu2system.vhd(8[13:16])
    wire we_N_63 /* synthesis is_clock=1, SET_AS_NETWORK=\CPU/we_N_63 */ ;   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(13[13:15])
    wire [5:0]adress_5__N_3;
    
    wire clk_c_enable_10;
    wire [8:0]akku_o_8__N_44;
    wire [5:0]pc;   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(23[15:17])
    
    wire clk_c_enable_15, n2254, n742, clk_c_enable_3;
    wire [8:0]akku_o_8__N_11;
    wire [2:0]states;   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(25[15:21])
    
    wire n2245, n2;
    wire [5:0]pc_5__N_30_c;
    wire [2:0]states_2__N_53;
    
    wire n2246, n2252;
    wire [7:0]akku_o_8__N_36;
    
    wire n2256, n1488, n1487, n1486, n1485, n1484;
    
    FD1S3AX adreg_i1 (.D(adress_5__N_3[0]), .CK(clk_c), .Q(\adrram[0] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(29[9] 73[16])
    defparam adreg_i1.GSR = "ENABLED";
    FD1P3AX akku_i1 (.D(akku_o_8__N_44[0]), .SP(clk_c_enable_10), .CK(clk_c), 
            .Q(akku_o_c_0)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(29[9] 73[16])
    defparam akku_i1.GSR = "ENABLED";
    FD1P3AX pc_i0_i0 (.D(pc_5__N_30[0]), .SP(clk_c_enable_15), .CK(clk_c), 
            .Q(pc[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(29[9] 73[16])
    defparam pc_i0_i0.GSR = "ENABLED";
    LUT4 i664_2_lut_3_lut_4_lut (.A(data[7]), .B(akku_o_c_8), .C(n2254), 
         .D(data[6]), .Z(n742)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;
    defparam i664_2_lut_3_lut_4_lut.init = 16'hf8f0;
    FD1P3AX akku_i9 (.D(akku_o_8__N_11[8]), .SP(clk_c_enable_3), .CK(clk_c), 
            .Q(akku_o_c_8)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(29[9] 73[16])
    defparam akku_i9.GSR = "ENABLED";
    FD1P3AX akku_i8 (.D(akku_o_8__N_44[7]), .SP(clk_c_enable_10), .CK(clk_c), 
            .Q(akku_o_c_7)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(29[9] 73[16])
    defparam akku_i8.GSR = "ENABLED";
    FD1P3AX akku_i7 (.D(akku_o_8__N_44[6]), .SP(clk_c_enable_10), .CK(clk_c), 
            .Q(akku_o_c_6)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(29[9] 73[16])
    defparam akku_i7.GSR = "ENABLED";
    FD1P3AX akku_i6 (.D(akku_o_8__N_44[5]), .SP(clk_c_enable_10), .CK(clk_c), 
            .Q(akku_o_c_5)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(29[9] 73[16])
    defparam akku_i6.GSR = "ENABLED";
    FD1P3AX akku_i5 (.D(akku_o_8__N_44[4]), .SP(clk_c_enable_10), .CK(clk_c), 
            .Q(akku_o_c_4)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(29[9] 73[16])
    defparam akku_i5.GSR = "ENABLED";
    FD1P3AX akku_i4 (.D(akku_o_8__N_44[3]), .SP(clk_c_enable_10), .CK(clk_c), 
            .Q(akku_o_c_3)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(29[9] 73[16])
    defparam akku_i4.GSR = "ENABLED";
    FD1P3AX akku_i3 (.D(akku_o_8__N_44[2]), .SP(clk_c_enable_10), .CK(clk_c), 
            .Q(akku_o_c_2)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(29[9] 73[16])
    defparam akku_i3.GSR = "ENABLED";
    FD1S3IX states__i2 (.D(n2245), .CK(clk_c), .CD(n2254), .Q(states[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(29[9] 73[16])
    defparam states__i2.GSR = "ENABLED";
    FD1P3AX akku_i2 (.D(akku_o_8__N_44[1]), .SP(clk_c_enable_10), .CK(clk_c), 
            .Q(akku_o_c_1)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(29[9] 73[16])
    defparam akku_i2.GSR = "ENABLED";
    FD1S3AX adreg_i6 (.D(adress_5__N_3[5]), .CK(clk_c), .Q(\adrram[5] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(29[9] 73[16])
    defparam adreg_i6.GSR = "ENABLED";
    FD1S3AX adreg_i5 (.D(adress_5__N_3[4]), .CK(clk_c), .Q(\adrram[4] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(29[9] 73[16])
    defparam adreg_i5.GSR = "ENABLED";
    FD1S3AX adreg_i4 (.D(adress_5__N_3[3]), .CK(clk_c), .Q(\adrram[3] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(29[9] 73[16])
    defparam adreg_i4.GSR = "ENABLED";
    FD1S3AX adreg_i3 (.D(adress_5__N_3[2]), .CK(clk_c), .Q(\adrram[2] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(29[9] 73[16])
    defparam adreg_i3.GSR = "ENABLED";
    FD1S3AX adreg_i2 (.D(adress_5__N_3[1]), .CK(clk_c), .Q(\adrram[1] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(29[9] 73[16])
    defparam adreg_i2.GSR = "ENABLED";
    FD1S3IX states__i1 (.D(n2), .CK(clk_c), .CD(n742), .Q(states[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(29[9] 73[16])
    defparam states__i1.GSR = "ENABLED";
    FD1P3AX pc_i0_i5 (.D(pc_5__N_30_c[5]), .SP(clk_c_enable_15), .CK(clk_c), 
            .Q(pc[5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(29[9] 73[16])
    defparam pc_i0_i5.GSR = "ENABLED";
    FD1P3AX pc_i0_i4 (.D(pc_5__N_30_c[4]), .SP(clk_c_enable_15), .CK(clk_c), 
            .Q(pc[4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(29[9] 73[16])
    defparam pc_i0_i4.GSR = "ENABLED";
    FD1P3AX pc_i0_i3 (.D(pc_5__N_30_c[3]), .SP(clk_c_enable_15), .CK(clk_c), 
            .Q(pc[3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(29[9] 73[16])
    defparam pc_i0_i3.GSR = "ENABLED";
    FD1P3AX pc_i0_i2 (.D(pc_5__N_30_c[2]), .SP(clk_c_enable_15), .CK(clk_c), 
            .Q(pc[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(29[9] 73[16])
    defparam pc_i0_i2.GSR = "ENABLED";
    FD1P3AX pc_i0_i1 (.D(pc_5__N_30_c[1]), .SP(clk_c_enable_15), .CK(clk_c), 
            .Q(pc[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(29[9] 73[16])
    defparam pc_i0_i1.GSR = "ENABLED";
    FD1S3IX states__i0 (.D(states_2__N_53[0]), .CK(clk_c), .CD(n2254), 
            .Q(states[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(29[9] 73[16])
    defparam states__i0.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_15_3_lut (.A(data[7]), .B(akku_o_c_8), .C(data[6]), 
         .Z(n2245)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_rep_15_3_lut.init = 16'h8080;
    LUT4 pc_5__I_0_85_i1_3_lut (.A(data[0]), .B(pc[0]), .C(n2254), .Z(adress_5__N_3[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(37[13] 44[20])
    defparam pc_5__I_0_85_i1_3_lut.init = 16'hcaca;
    LUT4 i435_3_lut_4_lut (.A(\adrram[3] ), .B(n2246), .C(\adrram[4] ), 
         .D(\adrram[5] ), .Z(pc_5__N_30_c[5])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // E:/Diamond/diamond/3.10_x64/ispfpga/vhdl_packages/numeric_std.vhd(1241[12:13])
    defparam i435_3_lut_4_lut.init = 16'h7f80;
    LUT4 i428_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2252), .C(\adrram[4] ), 
         .D(\adrram[3] ), .Z(pc_5__N_30_c[4])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // E:/Diamond/diamond/3.10_x64/ispfpga/vhdl_packages/numeric_std.vhd(1241[12:13])
    defparam i428_2_lut_3_lut_4_lut.init = 16'h78f0;
    LUT4 i1131_2_lut (.A(akku_o_8__N_44[8]), .B(states[2]), .Z(akku_o_8__N_11[8])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(47[13] 53[22])
    defparam i1131_2_lut.init = 16'h2222;
    LUT4 pc_5__I_0_85_i6_3_lut (.A(data[5]), .B(pc[5]), .C(n2254), .Z(adress_5__N_3[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(37[13] 44[20])
    defparam pc_5__I_0_85_i6_3_lut.init = 16'hcaca;
    LUT4 pc_5__I_0_85_i5_3_lut (.A(data[4]), .B(pc[4]), .C(n2254), .Z(adress_5__N_3[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(37[13] 44[20])
    defparam pc_5__I_0_85_i5_3_lut.init = 16'hcaca;
    LUT4 pc_5__I_0_85_i4_3_lut (.A(data[3]), .B(pc[3]), .C(n2254), .Z(adress_5__N_3[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(37[13] 44[20])
    defparam pc_5__I_0_85_i4_3_lut.init = 16'hcaca;
    LUT4 pc_5__I_0_85_i3_3_lut (.A(data[2]), .B(pc[2]), .C(n2254), .Z(adress_5__N_3[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(37[13] 44[20])
    defparam pc_5__I_0_85_i3_3_lut.init = 16'hcaca;
    LUT4 pc_5__I_0_85_i2_3_lut (.A(data[1]), .B(pc[1]), .C(n2254), .Z(adress_5__N_3[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(37[13] 44[20])
    defparam pc_5__I_0_85_i2_3_lut.init = 16'hcaca;
    LUT4 i486_1_lut (.A(data[7]), .Z(n2)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(59[20:43])
    defparam i486_1_lut.init = 16'h5555;
    LUT4 i407_2_lut (.A(\adrram[1] ), .B(\adrram[0] ), .Z(pc_5__N_30_c[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // E:/Diamond/diamond/3.10_x64/ispfpga/vhdl_packages/numeric_std.vhd(1241[12:13])
    defparam i407_2_lut.init = 16'h6666;
    LUT4 i2231_2_lut (.A(akku_o_c_6), .B(data[6]), .Z(akku_o_8__N_36[6])) /* synthesis lut_function=(!(A+(B))) */ ;   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(50[60:94])
    defparam i2231_2_lut.init = 16'h1111;
    LUT4 i2228_2_lut (.A(akku_o_c_7), .B(data[7]), .Z(akku_o_8__N_36[7])) /* synthesis lut_function=(!(A+(B))) */ ;   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(50[60:94])
    defparam i2228_2_lut.init = 16'h1111;
    LUT4 i2237_2_lut (.A(akku_o_c_4), .B(data[4]), .Z(akku_o_8__N_36[4])) /* synthesis lut_function=(!(A+(B))) */ ;   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(50[60:94])
    defparam i2237_2_lut.init = 16'h1111;
    LUT4 i2234_2_lut (.A(akku_o_c_5), .B(data[5]), .Z(akku_o_8__N_36[5])) /* synthesis lut_function=(!(A+(B))) */ ;   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(50[60:94])
    defparam i2234_2_lut.init = 16'h1111;
    LUT4 i2243_2_lut (.A(akku_o_c_2), .B(data[2]), .Z(akku_o_8__N_36[2])) /* synthesis lut_function=(!(A+(B))) */ ;   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(50[60:94])
    defparam i2243_2_lut.init = 16'h1111;
    LUT4 i2240_2_lut (.A(akku_o_c_3), .B(data[3]), .Z(akku_o_8__N_36[3])) /* synthesis lut_function=(!(A+(B))) */ ;   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(50[60:94])
    defparam i2240_2_lut.init = 16'h1111;
    LUT4 i2200_2_lut (.A(akku_o_c_0), .B(data[0]), .Z(akku_o_8__N_36[0])) /* synthesis lut_function=(!(A+(B))) */ ;   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(50[60:94])
    defparam i2200_2_lut.init = 16'h1111;
    LUT4 i2176_2_lut (.A(akku_o_c_1), .B(data[1]), .Z(akku_o_8__N_36[1])) /* synthesis lut_function=(!(A+(B))) */ ;   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(50[60:94])
    defparam i2176_2_lut.init = 16'h1111;
    LUT4 i409_2_lut_rep_22 (.A(\adrram[1] ), .B(\adrram[0] ), .Z(n2252)) /* synthesis lut_function=(A (B)) */ ;   // E:/Diamond/diamond/3.10_x64/ispfpga/vhdl_packages/numeric_std.vhd(1241[12:13])
    defparam i409_2_lut_rep_22.init = 16'h8888;
    LUT4 i416_2_lut_rep_16_3_lut (.A(\adrram[1] ), .B(\adrram[0] ), .C(\adrram[2] ), 
         .Z(n2246)) /* synthesis lut_function=(A (B (C))) */ ;   // E:/Diamond/diamond/3.10_x64/ispfpga/vhdl_packages/numeric_std.vhd(1241[12:13])
    defparam i416_2_lut_rep_16_3_lut.init = 16'h8080;
    LUT4 i414_2_lut_3_lut (.A(\adrram[1] ), .B(\adrram[0] ), .C(\adrram[2] ), 
         .Z(pc_5__N_30_c[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // E:/Diamond/diamond/3.10_x64/ispfpga/vhdl_packages/numeric_std.vhd(1241[12:13])
    defparam i414_2_lut_3_lut.init = 16'h7878;
    LUT4 i421_2_lut_3_lut_4_lut (.A(\adrram[1] ), .B(\adrram[0] ), .C(\adrram[3] ), 
         .D(\adrram[2] ), .Z(pc_5__N_30_c[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // E:/Diamond/diamond/3.10_x64/ispfpga/vhdl_packages/numeric_std.vhd(1241[12:13])
    defparam i421_2_lut_3_lut_4_lut.init = 16'h78f0;
    LUT4 i671_2_lut_rep_23 (.A(states[1]), .B(states[2]), .Z(clk_c_enable_10)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(47[13] 53[22])
    defparam i671_2_lut_rep_23.init = 16'h2222;
    LUT4 i13_4_lut_3_lut (.A(states[1]), .B(states[2]), .C(states[0]), 
         .Z(clk_c_enable_3)) /* synthesis lut_function=(!(A (B+(C))+!A !(B (C)))) */ ;   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(47[13] 53[22])
    defparam i13_4_lut_3_lut.init = 16'h4242;
    LUT4 i2_3_lut_rep_24 (.A(states[2]), .B(states[0]), .C(states[1]), 
         .Z(n2254)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(56[17:32])
    defparam i2_3_lut_rep_24.init = 16'hfefe;
    LUT4 i800_1_lut_3_lut (.A(states[2]), .B(states[0]), .C(states[1]), 
         .Z(clk_c_enable_15)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(56[17:32])
    defparam i800_1_lut_3_lut.init = 16'h0101;
    LUT4 i1_2_lut_3_lut_4_lut (.A(reset_c), .B(clk_c), .C(n2256), .D(states[2]), 
         .Z(we_N_63)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(84[21:60])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0002;
    LUT4 i1_2_lut_rep_26 (.A(states[1]), .B(states[0]), .Z(n2256)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(84[21:60])
    defparam i1_2_lut_rep_26.init = 16'hbbbb;
    LUT4 i1_2_lut_rep_17_3_lut (.A(states[1]), .B(states[0]), .C(states[2]), 
         .Z(n2247)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(84[21:60])
    defparam i1_2_lut_rep_17_3_lut.init = 16'hfbfb;
    LUT4 i1_2_lut_3_lut_4_lut_adj_8 (.A(states[1]), .B(states[0]), .C(clk_c), 
         .D(reset_c), .Z(oe_N_57)) /* synthesis lut_function=(!(A (C+!(D))+!A (B+(C+!(D))))) */ ;   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(84[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_8.init = 16'h0b00;
    LUT4 i1126_2_lut_3_lut (.A(data[7]), .B(akku_o_c_8), .C(data[6]), 
         .Z(states_2__N_53[0])) /* synthesis lut_function=(A (B+!(C))+!A !(C)) */ ;
    defparam i1126_2_lut_3_lut.init = 16'h8f8f;
    CCU2D add_91_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n1488), 
          .S0(akku_o_8__N_44[8]));   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(48[39:69])
    defparam add_91_cout.INIT0 = 16'h0000;
    defparam add_91_cout.INIT1 = 16'h0000;
    defparam add_91_cout.INJECT1_0 = "NO";
    defparam add_91_cout.INJECT1_1 = "NO";
    CCU2D add_91_9 (.A0(data[6]), .B0(states[0]), .C0(akku_o_8__N_36[6]), 
          .D0(akku_o_c_6), .A1(data[7]), .B1(states[0]), .C1(akku_o_8__N_36[7]), 
          .D1(akku_o_c_7), .CIN(n1487), .COUT(n1488), .S0(akku_o_8__N_44[6]), 
          .S1(akku_o_8__N_44[7]));   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(48[39:69])
    defparam add_91_9.INIT0 = 16'hd1e2;
    defparam add_91_9.INIT1 = 16'hd1e2;
    defparam add_91_9.INJECT1_0 = "NO";
    defparam add_91_9.INJECT1_1 = "NO";
    CCU2D add_91_7 (.A0(data[4]), .B0(states[0]), .C0(akku_o_8__N_36[4]), 
          .D0(akku_o_c_4), .A1(data[5]), .B1(states[0]), .C1(akku_o_8__N_36[5]), 
          .D1(akku_o_c_5), .CIN(n1486), .COUT(n1487), .S0(akku_o_8__N_44[4]), 
          .S1(akku_o_8__N_44[5]));   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(48[39:69])
    defparam add_91_7.INIT0 = 16'hd1e2;
    defparam add_91_7.INIT1 = 16'hd1e2;
    defparam add_91_7.INJECT1_0 = "NO";
    defparam add_91_7.INJECT1_1 = "NO";
    CCU2D add_91_5 (.A0(data[2]), .B0(states[0]), .C0(akku_o_8__N_36[2]), 
          .D0(akku_o_c_2), .A1(data[3]), .B1(states[0]), .C1(akku_o_8__N_36[3]), 
          .D1(akku_o_c_3), .CIN(n1485), .COUT(n1486), .S0(akku_o_8__N_44[2]), 
          .S1(akku_o_8__N_44[3]));   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(48[39:69])
    defparam add_91_5.INIT0 = 16'hd1e2;
    defparam add_91_5.INIT1 = 16'hd1e2;
    defparam add_91_5.INJECT1_0 = "NO";
    defparam add_91_5.INJECT1_1 = "NO";
    CCU2D add_91_3 (.A0(data[0]), .B0(states[0]), .C0(akku_o_8__N_36[0]), 
          .D0(akku_o_c_0), .A1(data[1]), .B1(states[0]), .C1(akku_o_8__N_36[1]), 
          .D1(akku_o_c_1), .CIN(n1484), .COUT(n1485), .S0(akku_o_8__N_44[0]), 
          .S1(akku_o_8__N_44[1]));   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(48[39:69])
    defparam add_91_3.INIT0 = 16'hd1e2;
    defparam add_91_3.INIT1 = 16'hd1e2;
    defparam add_91_3.INJECT1_0 = "NO";
    defparam add_91_3.INJECT1_1 = "NO";
    CCU2D add_91_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(states[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n1484));   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(48[39:69])
    defparam add_91_1.INIT0 = 16'hF000;
    defparam add_91_1.INIT1 = 16'h0fff;
    defparam add_91_1.INJECT1_0 = "NO";
    defparam add_91_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module TSALL
// module not written out since it is a black-box. 
//

//
// Verilog Description of module sram64kx8
//

module sram64kx8 (we_N_63, data, \adrram[5] , \adrram[3] , \adrram[2] , 
            \adrram[0] , akku_o_c_0, oe_N_57, n2247, akku_o_c_2, akku_o_c_7, 
            \adrram[1] , akku_o_c_6, \adrram[4] , \pc_5__N_30[0] , akku_o_c_1, 
            akku_o_c_5, akku_o_c_4, akku_o_c_3);
    input we_N_63;
    output [7:0]data;
    input \adrram[5] ;
    input \adrram[3] ;
    input \adrram[2] ;
    input \adrram[0] ;
    input akku_o_c_0;
    input oe_N_57;
    input n2247;
    input akku_o_c_2;
    input akku_o_c_7;
    input \adrram[1] ;
    input akku_o_c_6;
    input \adrram[4] ;
    output \pc_5__N_30[0] ;
    input akku_o_c_1;
    input akku_o_c_5;
    input akku_o_c_4;
    input akku_o_c_3;
    
    wire we_N_63 /* synthesis is_clock=1, SET_AS_NETWORK=\CPU/we_N_63 */ ;   // c:/users/70735/desktop/cpu_l/tb02cpu2.vhd(13[13:15])
    wire [7:0]\mem[22] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_414;
    wire [7:0]\mem[21] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_407;
    wire [7:0]\mem[53] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_512;
    wire [7:0]\mem[42] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_123;
    wire [7:0]\mem[52] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_133;
    wire [7:0]\mem[41] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_122;
    wire [7:0]\mem[40] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_121;
    wire [7:0]\mem[39] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_120;
    wire [7:0]\mem[23] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_376, n1783, n1814;
    wire [7:0]data_7__N_66;
    wire [7:0]\mem[38] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_119;
    wire [7:0]\mem[37] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_118;
    wire [7:0]\mem[36] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_117;
    wire [7:0]\mem[47] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_416;
    wire [7:0]\mem[35] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_107;
    wire [7:0]\mem[34] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_106;
    wire [7:0]\mem[51] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_373;
    wire [7:0]\mem[33] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_144;
    wire [7:0]\mem[2] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_168;
    wire [7:0]\mem[3] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_175;
    wire [7:0]\mem[4] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_182;
    wire [7:0]\mem[5] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_189;
    wire [7:0]\mem[6] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_196;
    wire [7:0]\mem[7] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_203;
    wire [7:0]\mem[8] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_210;
    wire [7:0]\mem[9] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_217;
    wire [7:0]\mem[10] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_224;
    wire [7:0]\mem[11] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_231;
    wire [7:0]\mem[12] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_238;
    wire [7:0]\mem[13] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_245;
    wire [7:0]\mem[14] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_252;
    wire [7:0]\mem[15] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_259;
    wire [7:0]\mem[16] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_266;
    wire [7:0]\mem[17] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_273;
    wire [7:0]\mem[18] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_280;
    wire [7:0]\mem[19] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_287;
    wire [7:0]\mem[20] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_294;
    wire [7:0]\mem[24] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_301;
    wire [7:0]\mem[25] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_308;
    wire [7:0]\mem[26] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_315;
    wire [7:0]\mem[27] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_322;
    wire [7:0]\mem[28] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_329;
    wire [7:0]\mem[29] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_336;
    wire [7:0]\mem[30] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_343;
    wire [7:0]\mem[31] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_350;
    wire [7:0]\mem[32] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_357;
    wire [7:0]\mem[63] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_364;
    wire [7:0]\mem[43] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_511;
    wire [7:0]\mem[44] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_475;
    wire [7:0]\mem[45] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_446;
    wire [7:0]\mem[46] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_423;
    wire [7:0]\mem[48] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_396;
    wire [7:0]\mem[49] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_389;
    wire [7:0]\mem[50] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_382;
    wire [7:0]\mem[54] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_505;
    wire [7:0]\mem[55] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_497;
    wire [7:0]\mem[56] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_488;
    wire [7:0]\mem[57] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_479;
    wire [7:0]\mem[58] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_470;
    wire [7:0]\mem[59] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_461;
    wire [7:0]\mem[60] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_452;
    wire [7:0]\mem[61] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_443;
    wire [7:0]\mem[62] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_433, n1752, n1845;
    wire [7:0]\mem[1] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_161;
    wire [7:0]\mem[0] ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(60[12:15])
    
    wire we_N_63_enable_154, n1721, n1876, n1690, n1907, n1659, 
        n1938, n1628, n1969, n1597, n2000, n1566, n2031, n1622, 
        n1623, n1626, n1624, n1625, n1627, n1686, n1687, n1689, 
        n1684, n1685, n1688, n1808, n1809, n1812, n1810, n1811, 
        n1813, n1932, n1933, n1936, n1934, n1935, n1937, n1994, 
        n1995, n1998, n1560, n1561, n1564, n1996, n1997, n1999, 
        n1839, n1840, n1843, n1841, n1842, n1844, n1591, n1592, 
        n1595, n1562, n1563, n1565, n1593, n1594, n1596, n2025, 
        n2026, n2029, n2027, n2028, n2030, n1653, n1654, n1657, 
        n1655, n1656, n1658, n1870, n1871, n1874, n1872, n1873, 
        n1875, n1963, n1964, n1967, n1965, n1966, n1968, n1715, 
        n1716, n1719, n1717, n1718, n1720, n1746, n1747, n1750, 
        n1748, n1749, n1751, n1901, n1902, n1905, n1903, n1904, 
        n1906, n1777, n1778, n1781, n1779, n1780, n1782, n1614, 
        n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1552, 
        n1553, n1554, n1555, n1556, n1557, n1800, n1801, n1924, 
        n1925, n1802, n1803, n1804, n1805, n1986, n1987, n1926, 
        n1927, n1568, n1806, n1807, n1682, n1683, n1928, n1929, 
        n1680, n1681, n1678, n1679, n1676, n1677, n2017, n2018, 
        n1988, n1989, n1930, n1931, n1990, n1991, n2019, n2020, 
        n1992, n1993, n1558, n1559, n1583, n1584, n1585, n1586, 
        n2021, n2022, n1831, n1832, n2023, n2024, n1833, n1834, 
        n1835, n1836, n1567, n1645, n1646, n1837, n1838, n1647, 
        n1648, n1587, n1588, n1649, n1650, n1589, n1590, n1651, 
        n1652, n1862, n1863, n1851, n1955, n1956, n1672, n1673, 
        n1864, n1865, n1866, n1867, n1957, n1958, n1868, n1869, 
        n1959, n1960, n1961, n1962, n1850, n1707, n1708, n1709, 
        n1710, n1711, n1712, n1713, n1714, n1738, n1739, n1740, 
        n1741, n1849, n1742, n1743, n1893, n1894, n1744, n1745, 
        n1848, n1895, n1896, n1897, n1898, n1948, n1899, n1900, 
        n1769, n1770, n1771, n1772, n1773, n1774, n1947, n1775, 
        n1776, n1598, n1599, n1847, n1600, n1601, n1602, n1603, 
        n1846, n1604, n1605, n1546, n1547, n1946, n2011, n2012, 
        n1976, n1977, n1945, n1606, n1607, n1608, n1609, n1944, 
        n1943, n1610, n1611, n1612, n1613, n1545, n1544, n1908, 
        n1909, n1978, n1979, n1942, n1941, n1910, n1911, n1940, 
        n1939, n1543, n1542, n1541, n1540, n1912, n1913, n2013, 
        n2014, n1644, n1980, n1981, n1643, n1914, n1915, n1642, 
        n1641, n1784, n1785, n1640, n1639, n1916, n1917, n1638, 
        n1786, n1787, n1637, n1636, n1788, n1789, n1982, n1983, 
        n1635, n1579, n1580, n1634, n1581, n1582, n1633, n1830, 
        n1815, n1816, n1829, n1817, n1818, n1819, n1820, n1632, 
        n1631, n1949, n1950, n1539, n2008, n1573, n1574, n1538, 
        n1730, n1852, n1853, n2007, n1660, n1661, n2004, n1729, 
        n1569, n1570, n1971, n1951, n1952, n2003, n1571, n1572, 
        n1728, n1856, n1857, n1880, n1698, n2250, n2249, n1821, 
        n1822, n1970, n1879, n1537, n1886, n1697, n1666, n1768, 
        n1536, n1885, n1878, n1767, n1877, n1696, n1860, n1551, 
        n1727, n1695, n1665, n1855, n2248, n1766, n1550, n1726, 
        n1706, n1664, n1954, n1765, n1705, n1694, n1953, n1854, 
        n2002, n1764, n2001, n1725, n1763, n1892, n1724, n1891, 
        n1762, n1761, n1737, n1760, n1736, n1884, n1823, n1824, 
        n1825, n1826, n1704, n1827, n1828, n1629, n1630, n1693, 
        n1575, n1576, n1858, n1859, n1668, n1669, n1699, n1700, 
        n1670, n1671, n1759, n1674, n1675, n1798, n1799, n1890, 
        n1922, n1923, n1984, n1985, n1548, n1549, n1883, n1703, 
        n1889, n1758, n1757, n1663, n1735, n1756, n1734, n1723, 
        n1702, n1692, n1755, n1733, n1722, n1974, n1975, n1701, 
        n1691, n1662, n1732, n1754, n1753, n1578, n1888, n2006, 
        n1887, n1882, n1577, n2005, n1731, n1881, n1918, n1919, 
        n1790, n1791, n1792, n1793, n1920, n1921, n1794, n1795, 
        n2257, n1796, n1797, n2015, n2016, n2010, n2259, n2009, 
        n2258, n2251, n2255, n1973, n1972, n1667, n1861;
    
    FD1P3AX mem_22__i0_i0 (.D(data[0]), .SP(we_N_63_enable_414), .CK(we_N_63), 
            .Q(\mem[22] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_22__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_21__i0_i0 (.D(data[0]), .SP(we_N_63_enable_407), .CK(we_N_63), 
            .Q(\mem[21] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_21__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_53__i0_i2 (.D(data[2]), .SP(we_N_63_enable_512), .CK(we_N_63), 
            .Q(\mem[53] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_53__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_42__i0_i7 (.D(data[7]), .SP(we_N_63_enable_123), .CK(we_N_63), 
            .Q(\mem[42] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_42__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_42__i0_i6 (.D(data[6]), .SP(we_N_63_enable_123), .CK(we_N_63), 
            .Q(\mem[42] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_42__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_53__i0_i1 (.D(data[1]), .SP(we_N_63_enable_512), .CK(we_N_63), 
            .Q(\mem[53] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_53__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_42__i0_i5 (.D(data[5]), .SP(we_N_63_enable_123), .CK(we_N_63), 
            .Q(\mem[42] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_42__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_42__i0_i4 (.D(data[4]), .SP(we_N_63_enable_123), .CK(we_N_63), 
            .Q(\mem[42] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_42__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_52__i0_i7 (.D(data[7]), .SP(we_N_63_enable_133), .CK(we_N_63), 
            .Q(\mem[52] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_52__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_42__i0_i3 (.D(data[3]), .SP(we_N_63_enable_123), .CK(we_N_63), 
            .Q(\mem[42] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_42__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_42__i0_i2 (.D(data[2]), .SP(we_N_63_enable_123), .CK(we_N_63), 
            .Q(\mem[42] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_42__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_52__i0_i6 (.D(data[6]), .SP(we_N_63_enable_133), .CK(we_N_63), 
            .Q(\mem[52] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_52__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_42__i0_i1 (.D(data[1]), .SP(we_N_63_enable_123), .CK(we_N_63), 
            .Q(\mem[42] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_42__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_52__i0_i5 (.D(data[5]), .SP(we_N_63_enable_133), .CK(we_N_63), 
            .Q(\mem[52] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_52__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_41__i0_i7 (.D(data[7]), .SP(we_N_63_enable_122), .CK(we_N_63), 
            .Q(\mem[41] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_41__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_41__i0_i6 (.D(data[6]), .SP(we_N_63_enable_122), .CK(we_N_63), 
            .Q(\mem[41] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_41__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_52__i0_i4 (.D(data[4]), .SP(we_N_63_enable_133), .CK(we_N_63), 
            .Q(\mem[52] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_52__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_41__i0_i5 (.D(data[5]), .SP(we_N_63_enable_122), .CK(we_N_63), 
            .Q(\mem[41] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_41__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_41__i0_i4 (.D(data[4]), .SP(we_N_63_enable_122), .CK(we_N_63), 
            .Q(\mem[41] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_41__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_41__i0_i3 (.D(data[3]), .SP(we_N_63_enable_122), .CK(we_N_63), 
            .Q(\mem[41] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_41__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_41__i0_i2 (.D(data[2]), .SP(we_N_63_enable_122), .CK(we_N_63), 
            .Q(\mem[41] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_41__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_41__i0_i1 (.D(data[1]), .SP(we_N_63_enable_122), .CK(we_N_63), 
            .Q(\mem[41] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_41__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_40__i0_i7 (.D(data[7]), .SP(we_N_63_enable_121), .CK(we_N_63), 
            .Q(\mem[40] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_40__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_40__i0_i6 (.D(data[6]), .SP(we_N_63_enable_121), .CK(we_N_63), 
            .Q(\mem[40] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_40__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_40__i0_i5 (.D(data[5]), .SP(we_N_63_enable_121), .CK(we_N_63), 
            .Q(\mem[40] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_40__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_40__i0_i4 (.D(data[4]), .SP(we_N_63_enable_121), .CK(we_N_63), 
            .Q(\mem[40] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_40__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_40__i0_i3 (.D(data[3]), .SP(we_N_63_enable_121), .CK(we_N_63), 
            .Q(\mem[40] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_40__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_40__i0_i2 (.D(data[2]), .SP(we_N_63_enable_121), .CK(we_N_63), 
            .Q(\mem[40] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_40__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_40__i0_i1 (.D(data[1]), .SP(we_N_63_enable_121), .CK(we_N_63), 
            .Q(\mem[40] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_40__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_39__i0_i7 (.D(data[7]), .SP(we_N_63_enable_120), .CK(we_N_63), 
            .Q(\mem[39] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_39__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_39__i0_i6 (.D(data[6]), .SP(we_N_63_enable_120), .CK(we_N_63), 
            .Q(\mem[39] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_39__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_39__i0_i5 (.D(data[5]), .SP(we_N_63_enable_120), .CK(we_N_63), 
            .Q(\mem[39] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_39__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_39__i0_i4 (.D(data[4]), .SP(we_N_63_enable_120), .CK(we_N_63), 
            .Q(\mem[39] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_39__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_39__i0_i3 (.D(data[3]), .SP(we_N_63_enable_120), .CK(we_N_63), 
            .Q(\mem[39] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_39__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_39__i0_i2 (.D(data[2]), .SP(we_N_63_enable_120), .CK(we_N_63), 
            .Q(\mem[39] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_39__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_39__i0_i1 (.D(data[1]), .SP(we_N_63_enable_120), .CK(we_N_63), 
            .Q(\mem[39] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_39__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_23__i0_i0 (.D(data[0]), .SP(we_N_63_enable_376), .CK(we_N_63), 
            .Q(\mem[23] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_23__i0_i0.GSR = "ENABLED";
    PFUMX i119332_i1 (.BLUT(n1783), .ALUT(n1814), .C0(\adrram[5] ), .Z(data_7__N_66[7]));
    FD1P3AX mem_38__i0_i7 (.D(data[7]), .SP(we_N_63_enable_119), .CK(we_N_63), 
            .Q(\mem[38] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_38__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_38__i0_i6 (.D(data[6]), .SP(we_N_63_enable_119), .CK(we_N_63), 
            .Q(\mem[38] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_38__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_38__i0_i5 (.D(data[5]), .SP(we_N_63_enable_119), .CK(we_N_63), 
            .Q(\mem[38] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_38__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_52__i0_i3 (.D(data[3]), .SP(we_N_63_enable_133), .CK(we_N_63), 
            .Q(\mem[52] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_52__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_52__i0_i2 (.D(data[2]), .SP(we_N_63_enable_133), .CK(we_N_63), 
            .Q(\mem[52] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_52__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_38__i0_i4 (.D(data[4]), .SP(we_N_63_enable_119), .CK(we_N_63), 
            .Q(\mem[38] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_38__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_38__i0_i3 (.D(data[3]), .SP(we_N_63_enable_119), .CK(we_N_63), 
            .Q(\mem[38] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_38__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_38__i0_i2 (.D(data[2]), .SP(we_N_63_enable_119), .CK(we_N_63), 
            .Q(\mem[38] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_38__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_38__i0_i1 (.D(data[1]), .SP(we_N_63_enable_119), .CK(we_N_63), 
            .Q(\mem[38] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_38__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_37__i0_i7 (.D(data[7]), .SP(we_N_63_enable_118), .CK(we_N_63), 
            .Q(\mem[37] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_37__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_37__i0_i6 (.D(data[6]), .SP(we_N_63_enable_118), .CK(we_N_63), 
            .Q(\mem[37] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_37__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_37__i0_i5 (.D(data[5]), .SP(we_N_63_enable_118), .CK(we_N_63), 
            .Q(\mem[37] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_37__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_37__i0_i4 (.D(data[4]), .SP(we_N_63_enable_118), .CK(we_N_63), 
            .Q(\mem[37] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_37__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_37__i0_i3 (.D(data[3]), .SP(we_N_63_enable_118), .CK(we_N_63), 
            .Q(\mem[37] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_37__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_37__i0_i2 (.D(data[2]), .SP(we_N_63_enable_118), .CK(we_N_63), 
            .Q(\mem[37] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_37__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_37__i0_i1 (.D(data[1]), .SP(we_N_63_enable_118), .CK(we_N_63), 
            .Q(\mem[37] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_37__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_36__i0_i7 (.D(data[7]), .SP(we_N_63_enable_117), .CK(we_N_63), 
            .Q(\mem[36] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_36__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_36__i0_i6 (.D(data[6]), .SP(we_N_63_enable_117), .CK(we_N_63), 
            .Q(\mem[36] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_36__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_36__i0_i5 (.D(data[5]), .SP(we_N_63_enable_117), .CK(we_N_63), 
            .Q(\mem[36] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_36__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_36__i0_i4 (.D(data[4]), .SP(we_N_63_enable_117), .CK(we_N_63), 
            .Q(\mem[36] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_36__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_52__i0_i1 (.D(data[1]), .SP(we_N_63_enable_133), .CK(we_N_63), 
            .Q(\mem[52] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_52__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_36__i0_i3 (.D(data[3]), .SP(we_N_63_enable_117), .CK(we_N_63), 
            .Q(\mem[36] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_36__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_36__i0_i2 (.D(data[2]), .SP(we_N_63_enable_117), .CK(we_N_63), 
            .Q(\mem[36] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_36__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_47__i0_i4 (.D(data[4]), .SP(we_N_63_enable_416), .CK(we_N_63), 
            .Q(\mem[47] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_47__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_36__i0_i1 (.D(data[1]), .SP(we_N_63_enable_117), .CK(we_N_63), 
            .Q(\mem[36] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_36__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_35__i0_i7 (.D(data[7]), .SP(we_N_63_enable_107), .CK(we_N_63), 
            .Q(\mem[35] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_35__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_35__i0_i6 (.D(data[6]), .SP(we_N_63_enable_107), .CK(we_N_63), 
            .Q(\mem[35] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_35__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_35__i0_i5 (.D(data[5]), .SP(we_N_63_enable_107), .CK(we_N_63), 
            .Q(\mem[35] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_35__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_35__i0_i4 (.D(data[4]), .SP(we_N_63_enable_107), .CK(we_N_63), 
            .Q(\mem[35] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_35__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_35__i0_i3 (.D(data[3]), .SP(we_N_63_enable_107), .CK(we_N_63), 
            .Q(\mem[35] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_35__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_35__i0_i2 (.D(data[2]), .SP(we_N_63_enable_107), .CK(we_N_63), 
            .Q(\mem[35] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_35__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_35__i0_i1 (.D(data[1]), .SP(we_N_63_enable_107), .CK(we_N_63), 
            .Q(\mem[35] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_35__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_34__i0_i7 (.D(data[7]), .SP(we_N_63_enable_106), .CK(we_N_63), 
            .Q(\mem[34] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_34__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_34__i0_i6 (.D(data[6]), .SP(we_N_63_enable_106), .CK(we_N_63), 
            .Q(\mem[34] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_34__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_34__i0_i5 (.D(data[5]), .SP(we_N_63_enable_106), .CK(we_N_63), 
            .Q(\mem[34] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_34__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_34__i0_i4 (.D(data[4]), .SP(we_N_63_enable_106), .CK(we_N_63), 
            .Q(\mem[34] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_34__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_34__i0_i3 (.D(data[3]), .SP(we_N_63_enable_106), .CK(we_N_63), 
            .Q(\mem[34] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_34__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_34__i0_i2 (.D(data[2]), .SP(we_N_63_enable_106), .CK(we_N_63), 
            .Q(\mem[34] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_34__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_51__i0_i7 (.D(data[7]), .SP(we_N_63_enable_373), .CK(we_N_63), 
            .Q(\mem[51] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_51__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_34__i0_i1 (.D(data[1]), .SP(we_N_63_enable_106), .CK(we_N_63), 
            .Q(\mem[34] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_34__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_33__i0_i7 (.D(data[7]), .SP(we_N_63_enable_144), .CK(we_N_63), 
            .Q(\mem[33] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_33__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_51__i0_i6 (.D(data[6]), .SP(we_N_63_enable_373), .CK(we_N_63), 
            .Q(\mem[51] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_51__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_33__i0_i6 (.D(data[6]), .SP(we_N_63_enable_144), .CK(we_N_63), 
            .Q(\mem[33] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_33__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_33__i0_i5 (.D(data[5]), .SP(we_N_63_enable_144), .CK(we_N_63), 
            .Q(\mem[33] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_33__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_33__i0_i4 (.D(data[4]), .SP(we_N_63_enable_144), .CK(we_N_63), 
            .Q(\mem[33] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_33__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_33__i0_i3 (.D(data[3]), .SP(we_N_63_enable_144), .CK(we_N_63), 
            .Q(\mem[33] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_33__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_33__i0_i2 (.D(data[2]), .SP(we_N_63_enable_144), .CK(we_N_63), 
            .Q(\mem[33] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_33__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_2__i0 (.D(data[0]), .SP(we_N_63_enable_168), .CK(we_N_63), 
            .Q(\mem[2] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_2__i0.GSR = "ENABLED";
    FD1P3AX mem_3__i0 (.D(data[0]), .SP(we_N_63_enable_175), .CK(we_N_63), 
            .Q(\mem[3] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_3__i0.GSR = "ENABLED";
    FD1P3AX mem_4__i0 (.D(data[0]), .SP(we_N_63_enable_182), .CK(we_N_63), 
            .Q(\mem[4] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_4__i0.GSR = "ENABLED";
    FD1P3AY mem_5__i0 (.D(data[0]), .SP(we_N_63_enable_189), .CK(we_N_63), 
            .Q(\mem[5] [0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_5__i0.GSR = "ENABLED";
    FD1P3AX mem_6__i0 (.D(data[0]), .SP(we_N_63_enable_196), .CK(we_N_63), 
            .Q(\mem[6] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_6__i0.GSR = "ENABLED";
    FD1P3AY mem_7__i0 (.D(data[0]), .SP(we_N_63_enable_203), .CK(we_N_63), 
            .Q(\mem[7] [0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_7__i0.GSR = "ENABLED";
    FD1P3AY mem_8__i0 (.D(data[0]), .SP(we_N_63_enable_210), .CK(we_N_63), 
            .Q(\mem[8] [0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_8__i0.GSR = "ENABLED";
    FD1P3AX mem_9__i0 (.D(data[0]), .SP(we_N_63_enable_217), .CK(we_N_63), 
            .Q(\mem[9] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_9__i0.GSR = "ENABLED";
    FD1P3AX mem_10__i0 (.D(data[0]), .SP(we_N_63_enable_224), .CK(we_N_63), 
            .Q(\mem[10] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_10__i0.GSR = "ENABLED";
    FD1P3AX mem_11__i0 (.D(data[0]), .SP(we_N_63_enable_231), .CK(we_N_63), 
            .Q(\mem[11] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_11__i0.GSR = "ENABLED";
    FD1P3AX mem_12__i0 (.D(data[0]), .SP(we_N_63_enable_238), .CK(we_N_63), 
            .Q(\mem[12] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_12__i0.GSR = "ENABLED";
    FD1P3AX mem_13__i0 (.D(data[0]), .SP(we_N_63_enable_245), .CK(we_N_63), 
            .Q(\mem[13] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_13__i0.GSR = "ENABLED";
    FD1P3AY mem_14__i0 (.D(data[0]), .SP(we_N_63_enable_252), .CK(we_N_63), 
            .Q(\mem[14] [0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_14__i0.GSR = "ENABLED";
    FD1P3AX mem_15__i0 (.D(data[0]), .SP(we_N_63_enable_259), .CK(we_N_63), 
            .Q(\mem[15] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_15__i0.GSR = "ENABLED";
    FD1P3AY mem_16__i0 (.D(data[0]), .SP(we_N_63_enable_266), .CK(we_N_63), 
            .Q(\mem[16] [0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_16__i0.GSR = "ENABLED";
    FD1P3AX mem_17__i0 (.D(data[0]), .SP(we_N_63_enable_273), .CK(we_N_63), 
            .Q(\mem[17] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_17__i0.GSR = "ENABLED";
    FD1P3AX mem_18__i0 (.D(data[0]), .SP(we_N_63_enable_280), .CK(we_N_63), 
            .Q(\mem[18] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_18__i0.GSR = "ENABLED";
    FD1P3AY mem_19__i0 (.D(data[0]), .SP(we_N_63_enable_287), .CK(we_N_63), 
            .Q(\mem[19] [0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_19__i0.GSR = "ENABLED";
    FD1P3AY mem_20__i0 (.D(data[0]), .SP(we_N_63_enable_294), .CK(we_N_63), 
            .Q(\mem[20] [0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_20__i0.GSR = "ENABLED";
    FD1P3AX mem_24__i0 (.D(data[0]), .SP(we_N_63_enable_301), .CK(we_N_63), 
            .Q(\mem[24] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_24__i0.GSR = "ENABLED";
    FD1P3AX mem_33__i0_i0 (.D(data[0]), .SP(we_N_63_enable_144), .CK(we_N_63), 
            .Q(\mem[33] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_33__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_34__i0_i0 (.D(data[0]), .SP(we_N_63_enable_106), .CK(we_N_63), 
            .Q(\mem[34] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_34__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_35__i0_i0 (.D(data[0]), .SP(we_N_63_enable_107), .CK(we_N_63), 
            .Q(\mem[35] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_35__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_25__i0 (.D(data[0]), .SP(we_N_63_enable_308), .CK(we_N_63), 
            .Q(\mem[25] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_25__i0.GSR = "ENABLED";
    FD1P3AY mem_26__i0 (.D(data[0]), .SP(we_N_63_enable_315), .CK(we_N_63), 
            .Q(\mem[26] [0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_26__i0.GSR = "ENABLED";
    FD1P3AX mem_27__i0 (.D(data[0]), .SP(we_N_63_enable_322), .CK(we_N_63), 
            .Q(\mem[27] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_27__i0.GSR = "ENABLED";
    FD1P3AX mem_28__i0 (.D(data[0]), .SP(we_N_63_enable_329), .CK(we_N_63), 
            .Q(\mem[28] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_28__i0.GSR = "ENABLED";
    FD1P3AX mem_29__i0 (.D(data[0]), .SP(we_N_63_enable_336), .CK(we_N_63), 
            .Q(\mem[29] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_29__i0.GSR = "ENABLED";
    FD1P3AX mem_30__i0 (.D(data[0]), .SP(we_N_63_enable_343), .CK(we_N_63), 
            .Q(\mem[30] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_30__i0.GSR = "ENABLED";
    FD1P3AX mem_31__i0 (.D(data[0]), .SP(we_N_63_enable_350), .CK(we_N_63), 
            .Q(\mem[31] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_31__i0.GSR = "ENABLED";
    FD1P3AX mem_32__i0 (.D(data[0]), .SP(we_N_63_enable_357), .CK(we_N_63), 
            .Q(\mem[32] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_32__i0.GSR = "ENABLED";
    FD1P3AY mem_63__i0 (.D(data[0]), .SP(we_N_63_enable_364), .CK(we_N_63), 
            .Q(\mem[63] [0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_63__i0.GSR = "ENABLED";
    FD1P3AX mem_36__i0_i0 (.D(data[0]), .SP(we_N_63_enable_117), .CK(we_N_63), 
            .Q(\mem[36] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_36__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_37__i0_i0 (.D(data[0]), .SP(we_N_63_enable_118), .CK(we_N_63), 
            .Q(\mem[37] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_37__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_38__i0_i0 (.D(data[0]), .SP(we_N_63_enable_119), .CK(we_N_63), 
            .Q(\mem[38] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_38__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_39__i0_i0 (.D(data[0]), .SP(we_N_63_enable_120), .CK(we_N_63), 
            .Q(\mem[39] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_39__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_40__i0_i0 (.D(data[0]), .SP(we_N_63_enable_121), .CK(we_N_63), 
            .Q(\mem[40] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_40__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_41__i0_i0 (.D(data[0]), .SP(we_N_63_enable_122), .CK(we_N_63), 
            .Q(\mem[41] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_41__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_42__i0_i0 (.D(data[0]), .SP(we_N_63_enable_123), .CK(we_N_63), 
            .Q(\mem[42] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_42__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_43__i0_i0 (.D(data[0]), .SP(we_N_63_enable_511), .CK(we_N_63), 
            .Q(\mem[43] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_43__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_44__i0_i0 (.D(data[0]), .SP(we_N_63_enable_475), .CK(we_N_63), 
            .Q(\mem[44] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_44__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_45__i0_i0 (.D(data[0]), .SP(we_N_63_enable_446), .CK(we_N_63), 
            .Q(\mem[45] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_45__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_46__i0_i0 (.D(data[0]), .SP(we_N_63_enable_423), .CK(we_N_63), 
            .Q(\mem[46] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_46__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_47__i0_i0 (.D(data[0]), .SP(we_N_63_enable_416), .CK(we_N_63), 
            .Q(\mem[47] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_47__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_48__i0_i0 (.D(data[0]), .SP(we_N_63_enable_396), .CK(we_N_63), 
            .Q(\mem[48] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_48__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_49__i0_i0 (.D(data[0]), .SP(we_N_63_enable_389), .CK(we_N_63), 
            .Q(\mem[49] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_49__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_50__i0_i0 (.D(data[0]), .SP(we_N_63_enable_382), .CK(we_N_63), 
            .Q(\mem[50] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_50__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_51__i0_i0 (.D(data[0]), .SP(we_N_63_enable_373), .CK(we_N_63), 
            .Q(\mem[51] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_51__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_52__i0_i0 (.D(data[0]), .SP(we_N_63_enable_133), .CK(we_N_63), 
            .Q(\mem[52] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_52__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_53__i0_i0 (.D(data[0]), .SP(we_N_63_enable_512), .CK(we_N_63), 
            .Q(\mem[53] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_53__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_54__i0_i0 (.D(data[0]), .SP(we_N_63_enable_505), .CK(we_N_63), 
            .Q(\mem[54] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_54__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_55__i0_i0 (.D(data[0]), .SP(we_N_63_enable_497), .CK(we_N_63), 
            .Q(\mem[55] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_55__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_56__i0_i0 (.D(data[0]), .SP(we_N_63_enable_488), .CK(we_N_63), 
            .Q(\mem[56] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_56__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_57__i0_i0 (.D(data[0]), .SP(we_N_63_enable_479), .CK(we_N_63), 
            .Q(\mem[57] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_57__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_58__i0_i0 (.D(data[0]), .SP(we_N_63_enable_470), .CK(we_N_63), 
            .Q(\mem[58] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_58__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_59__i0_i0 (.D(data[0]), .SP(we_N_63_enable_461), .CK(we_N_63), 
            .Q(\mem[59] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_59__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_60__i0_i0 (.D(data[0]), .SP(we_N_63_enable_452), .CK(we_N_63), 
            .Q(\mem[60] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_60__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_61__i0_i0 (.D(data[0]), .SP(we_N_63_enable_443), .CK(we_N_63), 
            .Q(\mem[61] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_61__i0_i0.GSR = "ENABLED";
    FD1P3AY mem_62__i0_i0 (.D(data[0]), .SP(we_N_63_enable_433), .CK(we_N_63), 
            .Q(\mem[62] [0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_62__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_33__i0_i1 (.D(data[1]), .SP(we_N_63_enable_144), .CK(we_N_63), 
            .Q(\mem[33] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_33__i0_i1.GSR = "ENABLED";
    PFUMX i118729_i1 (.BLUT(n1752), .ALUT(n1845), .C0(\adrram[5] ), .Z(data_7__N_66[6]));
    FD1P3AX mem_23__i0_i7 (.D(data[7]), .SP(we_N_63_enable_376), .CK(we_N_63), 
            .Q(\mem[23] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_23__i0_i7.GSR = "ENABLED";
    FD1P3AY mem_1__i0 (.D(data[0]), .SP(we_N_63_enable_161), .CK(we_N_63), 
            .Q(\mem[1] [0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_1__i0.GSR = "ENABLED";
    FD1P3AX mem_0__i0 (.D(data[0]), .SP(we_N_63_enable_154), .CK(we_N_63), 
            .Q(\mem[0] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_0__i0.GSR = "ENABLED";
    FD1P3AY mem_0__i1 (.D(data[1]), .SP(we_N_63_enable_154), .CK(we_N_63), 
            .Q(\mem[0] [1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_0__i1.GSR = "ENABLED";
    FD1P3AY mem_0__i2 (.D(data[2]), .SP(we_N_63_enable_154), .CK(we_N_63), 
            .Q(\mem[0] [2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_0__i2.GSR = "ENABLED";
    FD1P3AY mem_0__i3 (.D(data[3]), .SP(we_N_63_enable_154), .CK(we_N_63), 
            .Q(\mem[0] [3])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_0__i3.GSR = "ENABLED";
    FD1P3AY mem_0__i4 (.D(data[4]), .SP(we_N_63_enable_154), .CK(we_N_63), 
            .Q(\mem[0] [4])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_0__i4.GSR = "ENABLED";
    FD1P3AY mem_0__i5 (.D(data[5]), .SP(we_N_63_enable_154), .CK(we_N_63), 
            .Q(\mem[0] [5])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_0__i5.GSR = "ENABLED";
    FD1P3AX mem_0__i6 (.D(data[6]), .SP(we_N_63_enable_154), .CK(we_N_63), 
            .Q(\mem[0] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_0__i6.GSR = "ENABLED";
    FD1P3AX mem_0__i7 (.D(data[7]), .SP(we_N_63_enable_154), .CK(we_N_63), 
            .Q(\mem[0] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_0__i7.GSR = "ENABLED";
    FD1P3AY mem_1__i1 (.D(data[1]), .SP(we_N_63_enable_161), .CK(we_N_63), 
            .Q(\mem[1] [1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_1__i1.GSR = "ENABLED";
    FD1P3AX mem_1__i2 (.D(data[2]), .SP(we_N_63_enable_161), .CK(we_N_63), 
            .Q(\mem[1] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_1__i2.GSR = "ENABLED";
    FD1P3AX mem_1__i3 (.D(data[3]), .SP(we_N_63_enable_161), .CK(we_N_63), 
            .Q(\mem[1] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_1__i3.GSR = "ENABLED";
    FD1P3AY mem_1__i4 (.D(data[4]), .SP(we_N_63_enable_161), .CK(we_N_63), 
            .Q(\mem[1] [4])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_1__i4.GSR = "ENABLED";
    FD1P3AX mem_1__i5 (.D(data[5]), .SP(we_N_63_enable_161), .CK(we_N_63), 
            .Q(\mem[1] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_1__i5.GSR = "ENABLED";
    FD1P3AY mem_1__i6 (.D(data[6]), .SP(we_N_63_enable_161), .CK(we_N_63), 
            .Q(\mem[1] [6])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_1__i6.GSR = "ENABLED";
    FD1P3AX mem_1__i7 (.D(data[7]), .SP(we_N_63_enable_161), .CK(we_N_63), 
            .Q(\mem[1] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_1__i7.GSR = "ENABLED";
    FD1P3AY mem_2__i1 (.D(data[1]), .SP(we_N_63_enable_168), .CK(we_N_63), 
            .Q(\mem[2] [1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_2__i1.GSR = "ENABLED";
    FD1P3AY mem_2__i2 (.D(data[2]), .SP(we_N_63_enable_168), .CK(we_N_63), 
            .Q(\mem[2] [2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_2__i2.GSR = "ENABLED";
    FD1P3AX mem_2__i3 (.D(data[3]), .SP(we_N_63_enable_168), .CK(we_N_63), 
            .Q(\mem[2] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_2__i3.GSR = "ENABLED";
    FD1P3AY mem_2__i4 (.D(data[4]), .SP(we_N_63_enable_168), .CK(we_N_63), 
            .Q(\mem[2] [4])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_2__i4.GSR = "ENABLED";
    FD1P3AX mem_2__i5 (.D(data[5]), .SP(we_N_63_enable_168), .CK(we_N_63), 
            .Q(\mem[2] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_2__i5.GSR = "ENABLED";
    FD1P3AX mem_2__i6 (.D(data[6]), .SP(we_N_63_enable_168), .CK(we_N_63), 
            .Q(\mem[2] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_2__i6.GSR = "ENABLED";
    FD1P3AY mem_2__i7 (.D(data[7]), .SP(we_N_63_enable_168), .CK(we_N_63), 
            .Q(\mem[2] [7])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_2__i7.GSR = "ENABLED";
    FD1P3AY mem_3__i1 (.D(data[1]), .SP(we_N_63_enable_175), .CK(we_N_63), 
            .Q(\mem[3] [1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_3__i1.GSR = "ENABLED";
    FD1P3AY mem_3__i2 (.D(data[2]), .SP(we_N_63_enable_175), .CK(we_N_63), 
            .Q(\mem[3] [2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_3__i2.GSR = "ENABLED";
    FD1P3AY mem_3__i3 (.D(data[3]), .SP(we_N_63_enable_175), .CK(we_N_63), 
            .Q(\mem[3] [3])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_3__i3.GSR = "ENABLED";
    FD1P3AY mem_3__i4 (.D(data[4]), .SP(we_N_63_enable_175), .CK(we_N_63), 
            .Q(\mem[3] [4])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_3__i4.GSR = "ENABLED";
    FD1P3AY mem_3__i5 (.D(data[5]), .SP(we_N_63_enable_175), .CK(we_N_63), 
            .Q(\mem[3] [5])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_3__i5.GSR = "ENABLED";
    FD1P3AX mem_3__i6 (.D(data[6]), .SP(we_N_63_enable_175), .CK(we_N_63), 
            .Q(\mem[3] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_3__i6.GSR = "ENABLED";
    FD1P3AX mem_3__i7 (.D(data[7]), .SP(we_N_63_enable_175), .CK(we_N_63), 
            .Q(\mem[3] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_3__i7.GSR = "ENABLED";
    FD1P3AX mem_4__i1 (.D(data[1]), .SP(we_N_63_enable_182), .CK(we_N_63), 
            .Q(\mem[4] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_4__i1.GSR = "ENABLED";
    FD1P3AY mem_4__i2 (.D(data[2]), .SP(we_N_63_enable_182), .CK(we_N_63), 
            .Q(\mem[4] [2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_4__i2.GSR = "ENABLED";
    FD1P3AX mem_4__i3 (.D(data[3]), .SP(we_N_63_enable_182), .CK(we_N_63), 
            .Q(\mem[4] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_4__i3.GSR = "ENABLED";
    FD1P3AY mem_4__i4 (.D(data[4]), .SP(we_N_63_enable_182), .CK(we_N_63), 
            .Q(\mem[4] [4])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_4__i4.GSR = "ENABLED";
    FD1P3AX mem_4__i5 (.D(data[5]), .SP(we_N_63_enable_182), .CK(we_N_63), 
            .Q(\mem[4] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_4__i5.GSR = "ENABLED";
    FD1P3AY mem_4__i6 (.D(data[6]), .SP(we_N_63_enable_182), .CK(we_N_63), 
            .Q(\mem[4] [6])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_4__i6.GSR = "ENABLED";
    FD1P3AX mem_4__i7 (.D(data[7]), .SP(we_N_63_enable_182), .CK(we_N_63), 
            .Q(\mem[4] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_4__i7.GSR = "ENABLED";
    FD1P3AY mem_5__i1 (.D(data[1]), .SP(we_N_63_enable_189), .CK(we_N_63), 
            .Q(\mem[5] [1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_5__i1.GSR = "ENABLED";
    FD1P3AY mem_5__i2 (.D(data[2]), .SP(we_N_63_enable_189), .CK(we_N_63), 
            .Q(\mem[5] [2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_5__i2.GSR = "ENABLED";
    FD1P3AX mem_5__i3 (.D(data[3]), .SP(we_N_63_enable_189), .CK(we_N_63), 
            .Q(\mem[5] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_5__i3.GSR = "ENABLED";
    FD1P3AY mem_5__i4 (.D(data[4]), .SP(we_N_63_enable_189), .CK(we_N_63), 
            .Q(\mem[5] [4])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_5__i4.GSR = "ENABLED";
    FD1P3AX mem_5__i5 (.D(data[5]), .SP(we_N_63_enable_189), .CK(we_N_63), 
            .Q(\mem[5] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_5__i5.GSR = "ENABLED";
    FD1P3AX mem_5__i6 (.D(data[6]), .SP(we_N_63_enable_189), .CK(we_N_63), 
            .Q(\mem[5] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_5__i6.GSR = "ENABLED";
    FD1P3AY mem_5__i7 (.D(data[7]), .SP(we_N_63_enable_189), .CK(we_N_63), 
            .Q(\mem[5] [7])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_5__i7.GSR = "ENABLED";
    FD1P3AY mem_6__i1 (.D(data[1]), .SP(we_N_63_enable_196), .CK(we_N_63), 
            .Q(\mem[6] [1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_6__i1.GSR = "ENABLED";
    FD1P3AY mem_6__i2 (.D(data[2]), .SP(we_N_63_enable_196), .CK(we_N_63), 
            .Q(\mem[6] [2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_6__i2.GSR = "ENABLED";
    FD1P3AY mem_6__i3 (.D(data[3]), .SP(we_N_63_enable_196), .CK(we_N_63), 
            .Q(\mem[6] [3])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_6__i3.GSR = "ENABLED";
    FD1P3AY mem_6__i4 (.D(data[4]), .SP(we_N_63_enable_196), .CK(we_N_63), 
            .Q(\mem[6] [4])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_6__i4.GSR = "ENABLED";
    FD1P3AY mem_6__i5 (.D(data[5]), .SP(we_N_63_enable_196), .CK(we_N_63), 
            .Q(\mem[6] [5])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_6__i5.GSR = "ENABLED";
    FD1P3AX mem_6__i6 (.D(data[6]), .SP(we_N_63_enable_196), .CK(we_N_63), 
            .Q(\mem[6] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_6__i6.GSR = "ENABLED";
    FD1P3AX mem_6__i7 (.D(data[7]), .SP(we_N_63_enable_196), .CK(we_N_63), 
            .Q(\mem[6] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_6__i7.GSR = "ENABLED";
    FD1P3AY mem_7__i1 (.D(data[1]), .SP(we_N_63_enable_203), .CK(we_N_63), 
            .Q(\mem[7] [1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_7__i1.GSR = "ENABLED";
    FD1P3AY mem_7__i2 (.D(data[2]), .SP(we_N_63_enable_203), .CK(we_N_63), 
            .Q(\mem[7] [2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_7__i2.GSR = "ENABLED";
    FD1P3AX mem_7__i3 (.D(data[3]), .SP(we_N_63_enable_203), .CK(we_N_63), 
            .Q(\mem[7] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_7__i3.GSR = "ENABLED";
    FD1P3AY mem_7__i4 (.D(data[4]), .SP(we_N_63_enable_203), .CK(we_N_63), 
            .Q(\mem[7] [4])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_7__i4.GSR = "ENABLED";
    FD1P3AX mem_7__i5 (.D(data[5]), .SP(we_N_63_enable_203), .CK(we_N_63), 
            .Q(\mem[7] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_7__i5.GSR = "ENABLED";
    FD1P3AX mem_7__i6 (.D(data[6]), .SP(we_N_63_enable_203), .CK(we_N_63), 
            .Q(\mem[7] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_7__i6.GSR = "ENABLED";
    FD1P3AX mem_7__i7 (.D(data[7]), .SP(we_N_63_enable_203), .CK(we_N_63), 
            .Q(\mem[7] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_7__i7.GSR = "ENABLED";
    FD1P3AY mem_8__i1 (.D(data[1]), .SP(we_N_63_enable_210), .CK(we_N_63), 
            .Q(\mem[8] [1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_8__i1.GSR = "ENABLED";
    FD1P3AY mem_8__i2 (.D(data[2]), .SP(we_N_63_enable_210), .CK(we_N_63), 
            .Q(\mem[8] [2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_8__i2.GSR = "ENABLED";
    FD1P3AY mem_8__i3 (.D(data[3]), .SP(we_N_63_enable_210), .CK(we_N_63), 
            .Q(\mem[8] [3])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_8__i3.GSR = "ENABLED";
    FD1P3AY mem_8__i4 (.D(data[4]), .SP(we_N_63_enable_210), .CK(we_N_63), 
            .Q(\mem[8] [4])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_8__i4.GSR = "ENABLED";
    FD1P3AY mem_8__i5 (.D(data[5]), .SP(we_N_63_enable_210), .CK(we_N_63), 
            .Q(\mem[8] [5])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_8__i5.GSR = "ENABLED";
    FD1P3AY mem_8__i6 (.D(data[6]), .SP(we_N_63_enable_210), .CK(we_N_63), 
            .Q(\mem[8] [6])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_8__i6.GSR = "ENABLED";
    FD1P3AX mem_8__i7 (.D(data[7]), .SP(we_N_63_enable_210), .CK(we_N_63), 
            .Q(\mem[8] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_8__i7.GSR = "ENABLED";
    FD1P3AY mem_9__i1 (.D(data[1]), .SP(we_N_63_enable_217), .CK(we_N_63), 
            .Q(\mem[9] [1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_9__i1.GSR = "ENABLED";
    FD1P3AY mem_9__i2 (.D(data[2]), .SP(we_N_63_enable_217), .CK(we_N_63), 
            .Q(\mem[9] [2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_9__i2.GSR = "ENABLED";
    FD1P3AX mem_9__i3 (.D(data[3]), .SP(we_N_63_enable_217), .CK(we_N_63), 
            .Q(\mem[9] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_9__i3.GSR = "ENABLED";
    FD1P3AY mem_9__i4 (.D(data[4]), .SP(we_N_63_enable_217), .CK(we_N_63), 
            .Q(\mem[9] [4])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_9__i4.GSR = "ENABLED";
    FD1P3AX mem_9__i5 (.D(data[5]), .SP(we_N_63_enable_217), .CK(we_N_63), 
            .Q(\mem[9] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_9__i5.GSR = "ENABLED";
    FD1P3AY mem_9__i6 (.D(data[6]), .SP(we_N_63_enable_217), .CK(we_N_63), 
            .Q(\mem[9] [6])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_9__i6.GSR = "ENABLED";
    FD1P3AX mem_9__i7 (.D(data[7]), .SP(we_N_63_enable_217), .CK(we_N_63), 
            .Q(\mem[9] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_9__i7.GSR = "ENABLED";
    FD1P3AX mem_10__i1 (.D(data[1]), .SP(we_N_63_enable_224), .CK(we_N_63), 
            .Q(\mem[10] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_10__i1.GSR = "ENABLED";
    FD1P3AX mem_10__i2 (.D(data[2]), .SP(we_N_63_enable_224), .CK(we_N_63), 
            .Q(\mem[10] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_10__i2.GSR = "ENABLED";
    FD1P3AY mem_10__i3 (.D(data[3]), .SP(we_N_63_enable_224), .CK(we_N_63), 
            .Q(\mem[10] [3])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_10__i3.GSR = "ENABLED";
    FD1P3AY mem_10__i4 (.D(data[4]), .SP(we_N_63_enable_224), .CK(we_N_63), 
            .Q(\mem[10] [4])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_10__i4.GSR = "ENABLED";
    FD1P3AX mem_10__i5 (.D(data[5]), .SP(we_N_63_enable_224), .CK(we_N_63), 
            .Q(\mem[10] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_10__i5.GSR = "ENABLED";
    FD1P3AY mem_10__i6 (.D(data[6]), .SP(we_N_63_enable_224), .CK(we_N_63), 
            .Q(\mem[10] [6])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_10__i6.GSR = "ENABLED";
    FD1P3AY mem_10__i7 (.D(data[7]), .SP(we_N_63_enable_224), .CK(we_N_63), 
            .Q(\mem[10] [7])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_10__i7.GSR = "ENABLED";
    FD1P3AY mem_11__i1 (.D(data[1]), .SP(we_N_63_enable_231), .CK(we_N_63), 
            .Q(\mem[11] [1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_11__i1.GSR = "ENABLED";
    FD1P3AY mem_11__i2 (.D(data[2]), .SP(we_N_63_enable_231), .CK(we_N_63), 
            .Q(\mem[11] [2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_11__i2.GSR = "ENABLED";
    FD1P3AY mem_11__i3 (.D(data[3]), .SP(we_N_63_enable_231), .CK(we_N_63), 
            .Q(\mem[11] [3])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_11__i3.GSR = "ENABLED";
    FD1P3AY mem_11__i4 (.D(data[4]), .SP(we_N_63_enable_231), .CK(we_N_63), 
            .Q(\mem[11] [4])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_11__i4.GSR = "ENABLED";
    FD1P3AY mem_11__i5 (.D(data[5]), .SP(we_N_63_enable_231), .CK(we_N_63), 
            .Q(\mem[11] [5])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_11__i5.GSR = "ENABLED";
    FD1P3AY mem_11__i6 (.D(data[6]), .SP(we_N_63_enable_231), .CK(we_N_63), 
            .Q(\mem[11] [6])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_11__i6.GSR = "ENABLED";
    FD1P3AX mem_11__i7 (.D(data[7]), .SP(we_N_63_enable_231), .CK(we_N_63), 
            .Q(\mem[11] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_11__i7.GSR = "ENABLED";
    FD1P3AY mem_12__i1 (.D(data[1]), .SP(we_N_63_enable_238), .CK(we_N_63), 
            .Q(\mem[12] [1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_12__i1.GSR = "ENABLED";
    FD1P3AY mem_12__i2 (.D(data[2]), .SP(we_N_63_enable_238), .CK(we_N_63), 
            .Q(\mem[12] [2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_12__i2.GSR = "ENABLED";
    FD1P3AY mem_12__i3 (.D(data[3]), .SP(we_N_63_enable_238), .CK(we_N_63), 
            .Q(\mem[12] [3])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_12__i3.GSR = "ENABLED";
    FD1P3AY mem_12__i4 (.D(data[4]), .SP(we_N_63_enable_238), .CK(we_N_63), 
            .Q(\mem[12] [4])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_12__i4.GSR = "ENABLED";
    FD1P3AX mem_12__i5 (.D(data[5]), .SP(we_N_63_enable_238), .CK(we_N_63), 
            .Q(\mem[12] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_12__i5.GSR = "ENABLED";
    FD1P3AY mem_12__i6 (.D(data[6]), .SP(we_N_63_enable_238), .CK(we_N_63), 
            .Q(\mem[12] [6])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_12__i6.GSR = "ENABLED";
    FD1P3AY mem_12__i7 (.D(data[7]), .SP(we_N_63_enable_238), .CK(we_N_63), 
            .Q(\mem[12] [7])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_12__i7.GSR = "ENABLED";
    FD1P3AY mem_13__i1 (.D(data[1]), .SP(we_N_63_enable_245), .CK(we_N_63), 
            .Q(\mem[13] [1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_13__i1.GSR = "ENABLED";
    FD1P3AY mem_13__i2 (.D(data[2]), .SP(we_N_63_enable_245), .CK(we_N_63), 
            .Q(\mem[13] [2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_13__i2.GSR = "ENABLED";
    FD1P3AY mem_13__i3 (.D(data[3]), .SP(we_N_63_enable_245), .CK(we_N_63), 
            .Q(\mem[13] [3])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_13__i3.GSR = "ENABLED";
    FD1P3AY mem_13__i4 (.D(data[4]), .SP(we_N_63_enable_245), .CK(we_N_63), 
            .Q(\mem[13] [4])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_13__i4.GSR = "ENABLED";
    FD1P3AY mem_13__i5 (.D(data[5]), .SP(we_N_63_enable_245), .CK(we_N_63), 
            .Q(\mem[13] [5])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_13__i5.GSR = "ENABLED";
    FD1P3AX mem_13__i6 (.D(data[6]), .SP(we_N_63_enable_245), .CK(we_N_63), 
            .Q(\mem[13] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_13__i6.GSR = "ENABLED";
    FD1P3AX mem_13__i7 (.D(data[7]), .SP(we_N_63_enable_245), .CK(we_N_63), 
            .Q(\mem[13] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_13__i7.GSR = "ENABLED";
    FD1P3AY mem_14__i1 (.D(data[1]), .SP(we_N_63_enable_252), .CK(we_N_63), 
            .Q(\mem[14] [1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_14__i1.GSR = "ENABLED";
    FD1P3AY mem_14__i2 (.D(data[2]), .SP(we_N_63_enable_252), .CK(we_N_63), 
            .Q(\mem[14] [2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_14__i2.GSR = "ENABLED";
    FD1P3AX mem_14__i3 (.D(data[3]), .SP(we_N_63_enable_252), .CK(we_N_63), 
            .Q(\mem[14] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_14__i3.GSR = "ENABLED";
    FD1P3AY mem_14__i4 (.D(data[4]), .SP(we_N_63_enable_252), .CK(we_N_63), 
            .Q(\mem[14] [4])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_14__i4.GSR = "ENABLED";
    FD1P3AX mem_14__i5 (.D(data[5]), .SP(we_N_63_enable_252), .CK(we_N_63), 
            .Q(\mem[14] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_14__i5.GSR = "ENABLED";
    FD1P3AY mem_14__i6 (.D(data[6]), .SP(we_N_63_enable_252), .CK(we_N_63), 
            .Q(\mem[14] [6])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_14__i6.GSR = "ENABLED";
    FD1P3AX mem_14__i7 (.D(data[7]), .SP(we_N_63_enable_252), .CK(we_N_63), 
            .Q(\mem[14] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_14__i7.GSR = "ENABLED";
    FD1P3AX mem_15__i1 (.D(data[1]), .SP(we_N_63_enable_259), .CK(we_N_63), 
            .Q(\mem[15] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_15__i1.GSR = "ENABLED";
    FD1P3AY mem_15__i2 (.D(data[2]), .SP(we_N_63_enable_259), .CK(we_N_63), 
            .Q(\mem[15] [2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_15__i2.GSR = "ENABLED";
    FD1P3AX mem_15__i3 (.D(data[3]), .SP(we_N_63_enable_259), .CK(we_N_63), 
            .Q(\mem[15] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_15__i3.GSR = "ENABLED";
    FD1P3AY mem_15__i4 (.D(data[4]), .SP(we_N_63_enable_259), .CK(we_N_63), 
            .Q(\mem[15] [4])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_15__i4.GSR = "ENABLED";
    FD1P3AX mem_15__i5 (.D(data[5]), .SP(we_N_63_enable_259), .CK(we_N_63), 
            .Q(\mem[15] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_15__i5.GSR = "ENABLED";
    FD1P3AY mem_15__i6 (.D(data[6]), .SP(we_N_63_enable_259), .CK(we_N_63), 
            .Q(\mem[15] [6])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_15__i6.GSR = "ENABLED";
    FD1P3AX mem_15__i7 (.D(data[7]), .SP(we_N_63_enable_259), .CK(we_N_63), 
            .Q(\mem[15] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_15__i7.GSR = "ENABLED";
    FD1P3AY mem_16__i1 (.D(data[1]), .SP(we_N_63_enable_266), .CK(we_N_63), 
            .Q(\mem[16] [1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_16__i1.GSR = "ENABLED";
    FD1P3AY mem_16__i2 (.D(data[2]), .SP(we_N_63_enable_266), .CK(we_N_63), 
            .Q(\mem[16] [2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_16__i2.GSR = "ENABLED";
    FD1P3AX mem_16__i3 (.D(data[3]), .SP(we_N_63_enable_266), .CK(we_N_63), 
            .Q(\mem[16] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_16__i3.GSR = "ENABLED";
    FD1P3AY mem_16__i4 (.D(data[4]), .SP(we_N_63_enable_266), .CK(we_N_63), 
            .Q(\mem[16] [4])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_16__i4.GSR = "ENABLED";
    FD1P3AX mem_16__i5 (.D(data[5]), .SP(we_N_63_enable_266), .CK(we_N_63), 
            .Q(\mem[16] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_16__i5.GSR = "ENABLED";
    FD1P3AX mem_16__i6 (.D(data[6]), .SP(we_N_63_enable_266), .CK(we_N_63), 
            .Q(\mem[16] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_16__i6.GSR = "ENABLED";
    FD1P3AY mem_16__i7 (.D(data[7]), .SP(we_N_63_enable_266), .CK(we_N_63), 
            .Q(\mem[16] [7])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_16__i7.GSR = "ENABLED";
    FD1P3AY mem_17__i1 (.D(data[1]), .SP(we_N_63_enable_273), .CK(we_N_63), 
            .Q(\mem[17] [1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_17__i1.GSR = "ENABLED";
    FD1P3AY mem_17__i2 (.D(data[2]), .SP(we_N_63_enable_273), .CK(we_N_63), 
            .Q(\mem[17] [2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_17__i2.GSR = "ENABLED";
    FD1P3AX mem_17__i3 (.D(data[3]), .SP(we_N_63_enable_273), .CK(we_N_63), 
            .Q(\mem[17] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_17__i3.GSR = "ENABLED";
    FD1P3AX mem_17__i4 (.D(data[4]), .SP(we_N_63_enable_273), .CK(we_N_63), 
            .Q(\mem[17] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_17__i4.GSR = "ENABLED";
    FD1P3AX mem_17__i5 (.D(data[5]), .SP(we_N_63_enable_273), .CK(we_N_63), 
            .Q(\mem[17] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_17__i5.GSR = "ENABLED";
    FD1P3AY mem_17__i6 (.D(data[6]), .SP(we_N_63_enable_273), .CK(we_N_63), 
            .Q(\mem[17] [6])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_17__i6.GSR = "ENABLED";
    FD1P3AY mem_17__i7 (.D(data[7]), .SP(we_N_63_enable_273), .CK(we_N_63), 
            .Q(\mem[17] [7])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_17__i7.GSR = "ENABLED";
    FD1P3AY mem_18__i1 (.D(data[1]), .SP(we_N_63_enable_280), .CK(we_N_63), 
            .Q(\mem[18] [1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_18__i1.GSR = "ENABLED";
    FD1P3AY mem_18__i2 (.D(data[2]), .SP(we_N_63_enable_280), .CK(we_N_63), 
            .Q(\mem[18] [2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_18__i2.GSR = "ENABLED";
    FD1P3AX mem_18__i3 (.D(data[3]), .SP(we_N_63_enable_280), .CK(we_N_63), 
            .Q(\mem[18] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_18__i3.GSR = "ENABLED";
    FD1P3AX mem_18__i4 (.D(data[4]), .SP(we_N_63_enable_280), .CK(we_N_63), 
            .Q(\mem[18] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_18__i4.GSR = "ENABLED";
    FD1P3AX mem_18__i5 (.D(data[5]), .SP(we_N_63_enable_280), .CK(we_N_63), 
            .Q(\mem[18] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_18__i5.GSR = "ENABLED";
    FD1P3AY mem_18__i6 (.D(data[6]), .SP(we_N_63_enable_280), .CK(we_N_63), 
            .Q(\mem[18] [6])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_18__i6.GSR = "ENABLED";
    FD1P3AY mem_18__i7 (.D(data[7]), .SP(we_N_63_enable_280), .CK(we_N_63), 
            .Q(\mem[18] [7])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_18__i7.GSR = "ENABLED";
    FD1P3AX mem_19__i1 (.D(data[1]), .SP(we_N_63_enable_287), .CK(we_N_63), 
            .Q(\mem[19] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_19__i1.GSR = "ENABLED";
    FD1P3AX mem_19__i2 (.D(data[2]), .SP(we_N_63_enable_287), .CK(we_N_63), 
            .Q(\mem[19] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_19__i2.GSR = "ENABLED";
    FD1P3AY mem_19__i3 (.D(data[3]), .SP(we_N_63_enable_287), .CK(we_N_63), 
            .Q(\mem[19] [3])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_19__i3.GSR = "ENABLED";
    FD1P3AX mem_19__i4 (.D(data[4]), .SP(we_N_63_enable_287), .CK(we_N_63), 
            .Q(\mem[19] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_19__i4.GSR = "ENABLED";
    FD1P3AX mem_19__i5 (.D(data[5]), .SP(we_N_63_enable_287), .CK(we_N_63), 
            .Q(\mem[19] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_19__i5.GSR = "ENABLED";
    FD1P3AX mem_19__i6 (.D(data[6]), .SP(we_N_63_enable_287), .CK(we_N_63), 
            .Q(\mem[19] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_19__i6.GSR = "ENABLED";
    FD1P3AX mem_19__i7 (.D(data[7]), .SP(we_N_63_enable_287), .CK(we_N_63), 
            .Q(\mem[19] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_19__i7.GSR = "ENABLED";
    FD1P3AY mem_20__i1 (.D(data[1]), .SP(we_N_63_enable_294), .CK(we_N_63), 
            .Q(\mem[20] [1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_20__i1.GSR = "ENABLED";
    FD1P3AY mem_20__i2 (.D(data[2]), .SP(we_N_63_enable_294), .CK(we_N_63), 
            .Q(\mem[20] [2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_20__i2.GSR = "ENABLED";
    FD1P3AY mem_20__i3 (.D(data[3]), .SP(we_N_63_enable_294), .CK(we_N_63), 
            .Q(\mem[20] [3])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_20__i3.GSR = "ENABLED";
    FD1P3AX mem_20__i4 (.D(data[4]), .SP(we_N_63_enable_294), .CK(we_N_63), 
            .Q(\mem[20] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_20__i4.GSR = "ENABLED";
    FD1P3AX mem_20__i5 (.D(data[5]), .SP(we_N_63_enable_294), .CK(we_N_63), 
            .Q(\mem[20] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_20__i5.GSR = "ENABLED";
    FD1P3AX mem_20__i6 (.D(data[6]), .SP(we_N_63_enable_294), .CK(we_N_63), 
            .Q(\mem[20] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_20__i6.GSR = "ENABLED";
    FD1P3AX mem_20__i7 (.D(data[7]), .SP(we_N_63_enable_294), .CK(we_N_63), 
            .Q(\mem[20] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_20__i7.GSR = "ENABLED";
    FD1P3AY mem_24__i1 (.D(data[1]), .SP(we_N_63_enable_301), .CK(we_N_63), 
            .Q(\mem[24] [1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_24__i1.GSR = "ENABLED";
    FD1P3AY mem_24__i2 (.D(data[2]), .SP(we_N_63_enable_301), .CK(we_N_63), 
            .Q(\mem[24] [2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_24__i2.GSR = "ENABLED";
    FD1P3AY mem_24__i3 (.D(data[3]), .SP(we_N_63_enable_301), .CK(we_N_63), 
            .Q(\mem[24] [3])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_24__i3.GSR = "ENABLED";
    FD1P3AY mem_24__i4 (.D(data[4]), .SP(we_N_63_enable_301), .CK(we_N_63), 
            .Q(\mem[24] [4])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_24__i4.GSR = "ENABLED";
    FD1P3AY mem_24__i5 (.D(data[5]), .SP(we_N_63_enable_301), .CK(we_N_63), 
            .Q(\mem[24] [5])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_24__i5.GSR = "ENABLED";
    FD1P3AX mem_24__i6 (.D(data[6]), .SP(we_N_63_enable_301), .CK(we_N_63), 
            .Q(\mem[24] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_24__i6.GSR = "ENABLED";
    FD1P3AX mem_24__i7 (.D(data[7]), .SP(we_N_63_enable_301), .CK(we_N_63), 
            .Q(\mem[24] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_24__i7.GSR = "ENABLED";
    FD1P3AY mem_25__i1 (.D(data[1]), .SP(we_N_63_enable_308), .CK(we_N_63), 
            .Q(\mem[25] [1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_25__i1.GSR = "ENABLED";
    FD1P3AY mem_25__i2 (.D(data[2]), .SP(we_N_63_enable_308), .CK(we_N_63), 
            .Q(\mem[25] [2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_25__i2.GSR = "ENABLED";
    FD1P3AX mem_25__i3 (.D(data[3]), .SP(we_N_63_enable_308), .CK(we_N_63), 
            .Q(\mem[25] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_25__i3.GSR = "ENABLED";
    FD1P3AY mem_25__i4 (.D(data[4]), .SP(we_N_63_enable_308), .CK(we_N_63), 
            .Q(\mem[25] [4])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_25__i4.GSR = "ENABLED";
    FD1P3AX mem_25__i5 (.D(data[5]), .SP(we_N_63_enable_308), .CK(we_N_63), 
            .Q(\mem[25] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_25__i5.GSR = "ENABLED";
    FD1P3AY mem_25__i6 (.D(data[6]), .SP(we_N_63_enable_308), .CK(we_N_63), 
            .Q(\mem[25] [6])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_25__i6.GSR = "ENABLED";
    FD1P3AX mem_25__i7 (.D(data[7]), .SP(we_N_63_enable_308), .CK(we_N_63), 
            .Q(\mem[25] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_25__i7.GSR = "ENABLED";
    FD1P3AY mem_26__i1 (.D(data[1]), .SP(we_N_63_enable_315), .CK(we_N_63), 
            .Q(\mem[26] [1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_26__i1.GSR = "ENABLED";
    FD1P3AX mem_26__i2 (.D(data[2]), .SP(we_N_63_enable_315), .CK(we_N_63), 
            .Q(\mem[26] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_26__i2.GSR = "ENABLED";
    FD1P3AX mem_26__i3 (.D(data[3]), .SP(we_N_63_enable_315), .CK(we_N_63), 
            .Q(\mem[26] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_26__i3.GSR = "ENABLED";
    FD1P3AY mem_26__i4 (.D(data[4]), .SP(we_N_63_enable_315), .CK(we_N_63), 
            .Q(\mem[26] [4])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_26__i4.GSR = "ENABLED";
    FD1P3AX mem_26__i5 (.D(data[5]), .SP(we_N_63_enable_315), .CK(we_N_63), 
            .Q(\mem[26] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_26__i5.GSR = "ENABLED";
    FD1P3AY mem_26__i6 (.D(data[6]), .SP(we_N_63_enable_315), .CK(we_N_63), 
            .Q(\mem[26] [6])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_26__i6.GSR = "ENABLED";
    FD1P3AX mem_26__i7 (.D(data[7]), .SP(we_N_63_enable_315), .CK(we_N_63), 
            .Q(\mem[26] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_26__i7.GSR = "ENABLED";
    FD1P3AY mem_27__i1 (.D(data[1]), .SP(we_N_63_enable_322), .CK(we_N_63), 
            .Q(\mem[27] [1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_27__i1.GSR = "ENABLED";
    FD1P3AY mem_27__i2 (.D(data[2]), .SP(we_N_63_enable_322), .CK(we_N_63), 
            .Q(\mem[27] [2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_27__i2.GSR = "ENABLED";
    FD1P3AX mem_27__i3 (.D(data[3]), .SP(we_N_63_enable_322), .CK(we_N_63), 
            .Q(\mem[27] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_27__i3.GSR = "ENABLED";
    FD1P3AY mem_27__i4 (.D(data[4]), .SP(we_N_63_enable_322), .CK(we_N_63), 
            .Q(\mem[27] [4])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_27__i4.GSR = "ENABLED";
    FD1P3AX mem_27__i5 (.D(data[5]), .SP(we_N_63_enable_322), .CK(we_N_63), 
            .Q(\mem[27] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_27__i5.GSR = "ENABLED";
    FD1P3AX mem_27__i6 (.D(data[6]), .SP(we_N_63_enable_322), .CK(we_N_63), 
            .Q(\mem[27] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_27__i6.GSR = "ENABLED";
    FD1P3AY mem_27__i7 (.D(data[7]), .SP(we_N_63_enable_322), .CK(we_N_63), 
            .Q(\mem[27] [7])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_27__i7.GSR = "ENABLED";
    FD1P3AY mem_28__i1 (.D(data[1]), .SP(we_N_63_enable_329), .CK(we_N_63), 
            .Q(\mem[28] [1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_28__i1.GSR = "ENABLED";
    FD1P3AY mem_28__i2 (.D(data[2]), .SP(we_N_63_enable_329), .CK(we_N_63), 
            .Q(\mem[28] [2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_28__i2.GSR = "ENABLED";
    FD1P3AX mem_28__i3 (.D(data[3]), .SP(we_N_63_enable_329), .CK(we_N_63), 
            .Q(\mem[28] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_28__i3.GSR = "ENABLED";
    FD1P3AX mem_28__i4 (.D(data[4]), .SP(we_N_63_enable_329), .CK(we_N_63), 
            .Q(\mem[28] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_28__i4.GSR = "ENABLED";
    FD1P3AX mem_28__i5 (.D(data[5]), .SP(we_N_63_enable_329), .CK(we_N_63), 
            .Q(\mem[28] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_28__i5.GSR = "ENABLED";
    FD1P3AY mem_28__i6 (.D(data[6]), .SP(we_N_63_enable_329), .CK(we_N_63), 
            .Q(\mem[28] [6])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_28__i6.GSR = "ENABLED";
    FD1P3AY mem_28__i7 (.D(data[7]), .SP(we_N_63_enable_329), .CK(we_N_63), 
            .Q(\mem[28] [7])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_28__i7.GSR = "ENABLED";
    FD1P3AY mem_29__i1 (.D(data[1]), .SP(we_N_63_enable_336), .CK(we_N_63), 
            .Q(\mem[29] [1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_29__i1.GSR = "ENABLED";
    FD1P3AY mem_29__i2 (.D(data[2]), .SP(we_N_63_enable_336), .CK(we_N_63), 
            .Q(\mem[29] [2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_29__i2.GSR = "ENABLED";
    FD1P3AX mem_29__i3 (.D(data[3]), .SP(we_N_63_enable_336), .CK(we_N_63), 
            .Q(\mem[29] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_29__i3.GSR = "ENABLED";
    FD1P3AX mem_29__i4 (.D(data[4]), .SP(we_N_63_enable_336), .CK(we_N_63), 
            .Q(\mem[29] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_29__i4.GSR = "ENABLED";
    FD1P3AX mem_29__i5 (.D(data[5]), .SP(we_N_63_enable_336), .CK(we_N_63), 
            .Q(\mem[29] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_29__i5.GSR = "ENABLED";
    FD1P3AY mem_29__i6 (.D(data[6]), .SP(we_N_63_enable_336), .CK(we_N_63), 
            .Q(\mem[29] [6])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_29__i6.GSR = "ENABLED";
    FD1P3AY mem_29__i7 (.D(data[7]), .SP(we_N_63_enable_336), .CK(we_N_63), 
            .Q(\mem[29] [7])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_29__i7.GSR = "ENABLED";
    FD1P3AY mem_30__i1 (.D(data[1]), .SP(we_N_63_enable_343), .CK(we_N_63), 
            .Q(\mem[30] [1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_30__i1.GSR = "ENABLED";
    FD1P3AY mem_30__i2 (.D(data[2]), .SP(we_N_63_enable_343), .CK(we_N_63), 
            .Q(\mem[30] [2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_30__i2.GSR = "ENABLED";
    FD1P3AY mem_30__i3 (.D(data[3]), .SP(we_N_63_enable_343), .CK(we_N_63), 
            .Q(\mem[30] [3])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_30__i3.GSR = "ENABLED";
    FD1P3AY mem_30__i4 (.D(data[4]), .SP(we_N_63_enable_343), .CK(we_N_63), 
            .Q(\mem[30] [4])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_30__i4.GSR = "ENABLED";
    FD1P3AY mem_30__i5 (.D(data[5]), .SP(we_N_63_enable_343), .CK(we_N_63), 
            .Q(\mem[30] [5])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_30__i5.GSR = "ENABLED";
    FD1P3AX mem_30__i6 (.D(data[6]), .SP(we_N_63_enable_343), .CK(we_N_63), 
            .Q(\mem[30] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_30__i6.GSR = "ENABLED";
    FD1P3AX mem_30__i7 (.D(data[7]), .SP(we_N_63_enable_343), .CK(we_N_63), 
            .Q(\mem[30] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_30__i7.GSR = "ENABLED";
    FD1P3AY mem_31__i1 (.D(data[1]), .SP(we_N_63_enable_350), .CK(we_N_63), 
            .Q(\mem[31] [1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_31__i1.GSR = "ENABLED";
    FD1P3AY mem_31__i2 (.D(data[2]), .SP(we_N_63_enable_350), .CK(we_N_63), 
            .Q(\mem[31] [2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_31__i2.GSR = "ENABLED";
    FD1P3AX mem_31__i3 (.D(data[3]), .SP(we_N_63_enable_350), .CK(we_N_63), 
            .Q(\mem[31] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_31__i3.GSR = "ENABLED";
    FD1P3AY mem_31__i4 (.D(data[4]), .SP(we_N_63_enable_350), .CK(we_N_63), 
            .Q(\mem[31] [4])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_31__i4.GSR = "ENABLED";
    FD1P3AX mem_31__i5 (.D(data[5]), .SP(we_N_63_enable_350), .CK(we_N_63), 
            .Q(\mem[31] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_31__i5.GSR = "ENABLED";
    FD1P3AY mem_31__i6 (.D(data[6]), .SP(we_N_63_enable_350), .CK(we_N_63), 
            .Q(\mem[31] [6])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_31__i6.GSR = "ENABLED";
    FD1P3AX mem_31__i7 (.D(data[7]), .SP(we_N_63_enable_350), .CK(we_N_63), 
            .Q(\mem[31] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_31__i7.GSR = "ENABLED";
    FD1P3AX mem_32__i1 (.D(data[1]), .SP(we_N_63_enable_357), .CK(we_N_63), 
            .Q(\mem[32] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_32__i1.GSR = "ENABLED";
    FD1P3AX mem_32__i2 (.D(data[2]), .SP(we_N_63_enable_357), .CK(we_N_63), 
            .Q(\mem[32] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_32__i2.GSR = "ENABLED";
    FD1P3AX mem_32__i3 (.D(data[3]), .SP(we_N_63_enable_357), .CK(we_N_63), 
            .Q(\mem[32] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_32__i3.GSR = "ENABLED";
    FD1P3AX mem_32__i4 (.D(data[4]), .SP(we_N_63_enable_357), .CK(we_N_63), 
            .Q(\mem[32] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_32__i4.GSR = "ENABLED";
    FD1P3AY mem_32__i5 (.D(data[5]), .SP(we_N_63_enable_357), .CK(we_N_63), 
            .Q(\mem[32] [5])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_32__i5.GSR = "ENABLED";
    FD1P3AY mem_32__i6 (.D(data[6]), .SP(we_N_63_enable_357), .CK(we_N_63), 
            .Q(\mem[32] [6])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_32__i6.GSR = "ENABLED";
    FD1P3AY mem_32__i7 (.D(data[7]), .SP(we_N_63_enable_357), .CK(we_N_63), 
            .Q(\mem[32] [7])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_32__i7.GSR = "ENABLED";
    FD1P3AX mem_63__i1 (.D(data[1]), .SP(we_N_63_enable_364), .CK(we_N_63), 
            .Q(\mem[63] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_63__i1.GSR = "ENABLED";
    FD1P3AX mem_63__i2 (.D(data[2]), .SP(we_N_63_enable_364), .CK(we_N_63), 
            .Q(\mem[63] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_63__i2.GSR = "ENABLED";
    FD1P3AX mem_63__i3 (.D(data[3]), .SP(we_N_63_enable_364), .CK(we_N_63), 
            .Q(\mem[63] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_63__i3.GSR = "ENABLED";
    FD1P3AX mem_63__i4 (.D(data[4]), .SP(we_N_63_enable_364), .CK(we_N_63), 
            .Q(\mem[63] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_63__i4.GSR = "ENABLED";
    FD1P3AX mem_63__i5 (.D(data[5]), .SP(we_N_63_enable_364), .CK(we_N_63), 
            .Q(\mem[63] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_63__i5.GSR = "ENABLED";
    FD1P3AX mem_63__i6 (.D(data[6]), .SP(we_N_63_enable_364), .CK(we_N_63), 
            .Q(\mem[63] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_63__i6.GSR = "ENABLED";
    FD1P3AX mem_63__i7 (.D(data[7]), .SP(we_N_63_enable_364), .CK(we_N_63), 
            .Q(\mem[63] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_63__i7.GSR = "ENABLED";
    FD1P3AX mem_51__i0_i5 (.D(data[5]), .SP(we_N_63_enable_373), .CK(we_N_63), 
            .Q(\mem[51] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_51__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_23__i0_i6 (.D(data[6]), .SP(we_N_63_enable_376), .CK(we_N_63), 
            .Q(\mem[23] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_23__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_51__i0_i4 (.D(data[4]), .SP(we_N_63_enable_373), .CK(we_N_63), 
            .Q(\mem[51] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_51__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_23__i0_i5 (.D(data[5]), .SP(we_N_63_enable_376), .CK(we_N_63), 
            .Q(\mem[23] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_23__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_51__i0_i3 (.D(data[3]), .SP(we_N_63_enable_373), .CK(we_N_63), 
            .Q(\mem[51] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_51__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_23__i0_i4 (.D(data[4]), .SP(we_N_63_enable_376), .CK(we_N_63), 
            .Q(\mem[23] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_23__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_51__i0_i2 (.D(data[2]), .SP(we_N_63_enable_373), .CK(we_N_63), 
            .Q(\mem[51] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_51__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_23__i0_i3 (.D(data[3]), .SP(we_N_63_enable_376), .CK(we_N_63), 
            .Q(\mem[23] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_23__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_51__i0_i1 (.D(data[1]), .SP(we_N_63_enable_373), .CK(we_N_63), 
            .Q(\mem[51] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_51__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_23__i0_i2 (.D(data[2]), .SP(we_N_63_enable_376), .CK(we_N_63), 
            .Q(\mem[23] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_23__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_50__i0_i7 (.D(data[7]), .SP(we_N_63_enable_382), .CK(we_N_63), 
            .Q(\mem[50] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_50__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_23__i0_i1 (.D(data[1]), .SP(we_N_63_enable_376), .CK(we_N_63), 
            .Q(\mem[23] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_23__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_50__i0_i6 (.D(data[6]), .SP(we_N_63_enable_382), .CK(we_N_63), 
            .Q(\mem[50] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_50__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_50__i0_i5 (.D(data[5]), .SP(we_N_63_enable_382), .CK(we_N_63), 
            .Q(\mem[50] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_50__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_50__i0_i4 (.D(data[4]), .SP(we_N_63_enable_382), .CK(we_N_63), 
            .Q(\mem[50] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_50__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_50__i0_i3 (.D(data[3]), .SP(we_N_63_enable_382), .CK(we_N_63), 
            .Q(\mem[50] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_50__i0_i3.GSR = "ENABLED";
    PFUMX i118126_i1 (.BLUT(n1721), .ALUT(n1876), .C0(\adrram[5] ), .Z(data_7__N_66[5]));
    FD1P3AX mem_50__i0_i2 (.D(data[2]), .SP(we_N_63_enable_382), .CK(we_N_63), 
            .Q(\mem[50] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_50__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_50__i0_i1 (.D(data[1]), .SP(we_N_63_enable_382), .CK(we_N_63), 
            .Q(\mem[50] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_50__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_49__i0_i7 (.D(data[7]), .SP(we_N_63_enable_389), .CK(we_N_63), 
            .Q(\mem[49] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_49__i0_i7.GSR = "ENABLED";
    PFUMX i117523_i1 (.BLUT(n1690), .ALUT(n1907), .C0(\adrram[5] ), .Z(data_7__N_66[4]));
    FD1P3AX mem_49__i0_i6 (.D(data[6]), .SP(we_N_63_enable_389), .CK(we_N_63), 
            .Q(\mem[49] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_49__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_49__i0_i5 (.D(data[5]), .SP(we_N_63_enable_389), .CK(we_N_63), 
            .Q(\mem[49] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_49__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_49__i0_i4 (.D(data[4]), .SP(we_N_63_enable_389), .CK(we_N_63), 
            .Q(\mem[49] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_49__i0_i4.GSR = "ENABLED";
    PFUMX i116920_i1 (.BLUT(n1659), .ALUT(n1938), .C0(\adrram[5] ), .Z(data_7__N_66[3]));
    FD1P3AX mem_49__i0_i3 (.D(data[3]), .SP(we_N_63_enable_389), .CK(we_N_63), 
            .Q(\mem[49] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_49__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_49__i0_i2 (.D(data[2]), .SP(we_N_63_enable_389), .CK(we_N_63), 
            .Q(\mem[49] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_49__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_49__i0_i1 (.D(data[1]), .SP(we_N_63_enable_389), .CK(we_N_63), 
            .Q(\mem[49] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_49__i0_i1.GSR = "ENABLED";
    PFUMX i116317_i1 (.BLUT(n1628), .ALUT(n1969), .C0(\adrram[5] ), .Z(data_7__N_66[2]));
    FD1P3AX mem_48__i0_i7 (.D(data[7]), .SP(we_N_63_enable_396), .CK(we_N_63), 
            .Q(\mem[48] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_48__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_48__i0_i6 (.D(data[6]), .SP(we_N_63_enable_396), .CK(we_N_63), 
            .Q(\mem[48] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_48__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_48__i0_i5 (.D(data[5]), .SP(we_N_63_enable_396), .CK(we_N_63), 
            .Q(\mem[48] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_48__i0_i5.GSR = "ENABLED";
    PFUMX i115714_i1 (.BLUT(n1597), .ALUT(n2000), .C0(\adrram[5] ), .Z(data_7__N_66[1]));
    FD1P3AX mem_48__i0_i4 (.D(data[4]), .SP(we_N_63_enable_396), .CK(we_N_63), 
            .Q(\mem[48] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_48__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_48__i0_i3 (.D(data[3]), .SP(we_N_63_enable_396), .CK(we_N_63), 
            .Q(\mem[48] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_48__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_48__i0_i2 (.D(data[2]), .SP(we_N_63_enable_396), .CK(we_N_63), 
            .Q(\mem[48] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_48__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_48__i0_i1 (.D(data[1]), .SP(we_N_63_enable_396), .CK(we_N_63), 
            .Q(\mem[48] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_48__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_47__i0_i7 (.D(data[7]), .SP(we_N_63_enable_416), .CK(we_N_63), 
            .Q(\mem[47] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_47__i0_i7.GSR = "ENABLED";
    PFUMX i115111_i1 (.BLUT(n1566), .ALUT(n2031), .C0(\adrram[5] ), .Z(data_7__N_66[0]));
    L6MUX21 i1523 (.D0(n1622), .D1(n1623), .SD(\adrram[3] ), .Z(n1626));
    L6MUX21 i1524 (.D0(n1624), .D1(n1625), .SD(\adrram[3] ), .Z(n1627));
    L6MUX21 i1586 (.D0(n1686), .D1(n1687), .SD(\adrram[3] ), .Z(n1689));
    L6MUX21 i1585 (.D0(n1684), .D1(n1685), .SD(\adrram[3] ), .Z(n1688));
    L6MUX21 i1709 (.D0(n1808), .D1(n1809), .SD(\adrram[3] ), .Z(n1812));
    L6MUX21 i1710 (.D0(n1810), .D1(n1811), .SD(\adrram[3] ), .Z(n1813));
    L6MUX21 i1833 (.D0(n1932), .D1(n1933), .SD(\adrram[3] ), .Z(n1936));
    L6MUX21 i1834 (.D0(n1934), .D1(n1935), .SD(\adrram[3] ), .Z(n1937));
    L6MUX21 i1895 (.D0(n1994), .D1(n1995), .SD(\adrram[3] ), .Z(n1998));
    L6MUX21 i1461 (.D0(n1560), .D1(n1561), .SD(\adrram[3] ), .Z(n1564));
    L6MUX21 i1896 (.D0(n1996), .D1(n1997), .SD(\adrram[3] ), .Z(n1999));
    FD1P3AX mem_47__i0_i6 (.D(data[6]), .SP(we_N_63_enable_416), .CK(we_N_63), 
            .Q(\mem[47] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_47__i0_i6.GSR = "ENABLED";
    L6MUX21 i1740 (.D0(n1839), .D1(n1840), .SD(\adrram[3] ), .Z(n1843));
    L6MUX21 i1741 (.D0(n1841), .D1(n1842), .SD(\adrram[3] ), .Z(n1844));
    L6MUX21 i1492 (.D0(n1591), .D1(n1592), .SD(\adrram[3] ), .Z(n1595));
    L6MUX21 i1462 (.D0(n1562), .D1(n1563), .SD(\adrram[3] ), .Z(n1565));
    L6MUX21 i1493 (.D0(n1593), .D1(n1594), .SD(\adrram[3] ), .Z(n1596));
    L6MUX21 i1926 (.D0(n2025), .D1(n2026), .SD(\adrram[3] ), .Z(n2029));
    L6MUX21 i1927 (.D0(n2027), .D1(n2028), .SD(\adrram[3] ), .Z(n2030));
    FD1P3AX mem_47__i0_i5 (.D(data[5]), .SP(we_N_63_enable_416), .CK(we_N_63), 
            .Q(\mem[47] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_47__i0_i5.GSR = "ENABLED";
    L6MUX21 i1554 (.D0(n1653), .D1(n1654), .SD(\adrram[3] ), .Z(n1657));
    FD1P3AX mem_47__i0_i3 (.D(data[3]), .SP(we_N_63_enable_416), .CK(we_N_63), 
            .Q(\mem[47] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_47__i0_i3.GSR = "ENABLED";
    L6MUX21 i1555 (.D0(n1655), .D1(n1656), .SD(\adrram[3] ), .Z(n1658));
    L6MUX21 i1771 (.D0(n1870), .D1(n1871), .SD(\adrram[3] ), .Z(n1874));
    L6MUX21 i1772 (.D0(n1872), .D1(n1873), .SD(\adrram[3] ), .Z(n1875));
    L6MUX21 i1864 (.D0(n1963), .D1(n1964), .SD(\adrram[3] ), .Z(n1967));
    L6MUX21 i1865 (.D0(n1965), .D1(n1966), .SD(\adrram[3] ), .Z(n1968));
    L6MUX21 i1616 (.D0(n1715), .D1(n1716), .SD(\adrram[3] ), .Z(n1719));
    L6MUX21 i1617 (.D0(n1717), .D1(n1718), .SD(\adrram[3] ), .Z(n1720));
    L6MUX21 i1647 (.D0(n1746), .D1(n1747), .SD(\adrram[3] ), .Z(n1750));
    FD1P3AX mem_21__i0_i7 (.D(data[7]), .SP(we_N_63_enable_407), .CK(we_N_63), 
            .Q(\mem[21] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_21__i0_i7.GSR = "ENABLED";
    L6MUX21 i1648 (.D0(n1748), .D1(n1749), .SD(\adrram[3] ), .Z(n1751));
    L6MUX21 i1802 (.D0(n1901), .D1(n1902), .SD(\adrram[3] ), .Z(n1905));
    L6MUX21 i1803 (.D0(n1903), .D1(n1904), .SD(\adrram[3] ), .Z(n1906));
    L6MUX21 i1678 (.D0(n1777), .D1(n1778), .SD(\adrram[3] ), .Z(n1781));
    L6MUX21 i1679 (.D0(n1779), .D1(n1780), .SD(\adrram[3] ), .Z(n1782));
    FD1P3AX mem_21__i0_i6 (.D(data[6]), .SP(we_N_63_enable_407), .CK(we_N_63), 
            .Q(\mem[21] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_21__i0_i6.GSR = "ENABLED";
    L6MUX21 i1519 (.D0(n1614), .D1(n1615), .SD(\adrram[2] ), .Z(n1622));
    L6MUX21 i1520 (.D0(n1616), .D1(n1617), .SD(\adrram[2] ), .Z(n1623));
    L6MUX21 i1521 (.D0(n1618), .D1(n1619), .SD(\adrram[2] ), .Z(n1624));
    L6MUX21 i1522 (.D0(n1620), .D1(n1621), .SD(\adrram[2] ), .Z(n1625));
    L6MUX21 i1457 (.D0(n1552), .D1(n1553), .SD(\adrram[2] ), .Z(n1560));
    L6MUX21 i1458 (.D0(n1554), .D1(n1555), .SD(\adrram[2] ), .Z(n1561));
    FD1P3AX mem_21__i0_i5 (.D(data[5]), .SP(we_N_63_enable_407), .CK(we_N_63), 
            .Q(\mem[21] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_21__i0_i5.GSR = "ENABLED";
    L6MUX21 i1459 (.D0(n1556), .D1(n1557), .SD(\adrram[2] ), .Z(n1562));
    L6MUX21 i1705 (.D0(n1800), .D1(n1801), .SD(\adrram[2] ), .Z(n1808));
    L6MUX21 i1829 (.D0(n1924), .D1(n1925), .SD(\adrram[2] ), .Z(n1932));
    L6MUX21 i1706 (.D0(n1802), .D1(n1803), .SD(\adrram[2] ), .Z(n1809));
    L6MUX21 i1707 (.D0(n1804), .D1(n1805), .SD(\adrram[2] ), .Z(n1810));
    L6MUX21 i1891 (.D0(n1986), .D1(n1987), .SD(\adrram[2] ), .Z(n1994));
    L6MUX21 i1830 (.D0(n1926), .D1(n1927), .SD(\adrram[2] ), .Z(n1933));
    LUT4 i1465_3_lut (.A(\mem[2] [1]), .B(\mem[3] [1]), .C(\adrram[0] ), 
         .Z(n1568)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1465_3_lut.init = 16'hcaca;
    FD1P3AX mem_21__i0_i4 (.D(data[4]), .SP(we_N_63_enable_407), .CK(we_N_63), 
            .Q(\mem[21] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_21__i0_i4.GSR = "ENABLED";
    L6MUX21 i1708 (.D0(n1806), .D1(n1807), .SD(\adrram[2] ), .Z(n1811));
    L6MUX21 i1584 (.D0(n1682), .D1(n1683), .SD(\adrram[2] ), .Z(n1687));
    L6MUX21 i1831 (.D0(n1928), .D1(n1929), .SD(\adrram[2] ), .Z(n1934));
    L6MUX21 i1583 (.D0(n1680), .D1(n1681), .SD(\adrram[2] ), .Z(n1686));
    L6MUX21 i1582 (.D0(n1678), .D1(n1679), .SD(\adrram[2] ), .Z(n1685));
    L6MUX21 i1581 (.D0(n1676), .D1(n1677), .SD(\adrram[2] ), .Z(n1684));
    LUT4 Select_644_i3_4_lut (.A(data_7__N_66[0]), .B(akku_o_c_0), .C(oe_N_57), 
         .D(n2247), .Z(data[0])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((D)+!B)) */ ;
    defparam Select_644_i3_4_lut.init = 16'ha0ec;
    LUT4 Select_642_i3_4_lut (.A(data_7__N_66[2]), .B(akku_o_c_2), .C(oe_N_57), 
         .D(n2247), .Z(data[2])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((D)+!B)) */ ;
    defparam Select_642_i3_4_lut.init = 16'ha0ec;
    FD1P3AX mem_21__i0_i3 (.D(data[3]), .SP(we_N_63_enable_407), .CK(we_N_63), 
            .Q(\mem[21] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_21__i0_i3.GSR = "ENABLED";
    L6MUX21 i1922 (.D0(n2017), .D1(n2018), .SD(\adrram[2] ), .Z(n2025));
    L6MUX21 i1892 (.D0(n1988), .D1(n1989), .SD(\adrram[2] ), .Z(n1995));
    L6MUX21 i1832 (.D0(n1930), .D1(n1931), .SD(\adrram[2] ), .Z(n1935));
    L6MUX21 i1893 (.D0(n1990), .D1(n1991), .SD(\adrram[2] ), .Z(n1996));
    L6MUX21 i1923 (.D0(n2019), .D1(n2020), .SD(\adrram[2] ), .Z(n2026));
    L6MUX21 i1894 (.D0(n1992), .D1(n1993), .SD(\adrram[2] ), .Z(n1997));
    L6MUX21 i1460 (.D0(n1558), .D1(n1559), .SD(\adrram[2] ), .Z(n1563));
    LUT4 Select_637_i3_4_lut (.A(data_7__N_66[7]), .B(akku_o_c_7), .C(oe_N_57), 
         .D(n2247), .Z(data[7])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((D)+!B)) */ ;
    defparam Select_637_i3_4_lut.init = 16'ha0ec;
    FD1P3AX mem_21__i0_i2 (.D(data[2]), .SP(we_N_63_enable_407), .CK(we_N_63), 
            .Q(\mem[21] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_21__i0_i2.GSR = "ENABLED";
    L6MUX21 i1488 (.D0(n1583), .D1(n1584), .SD(\adrram[2] ), .Z(n1591));
    L6MUX21 i1489 (.D0(n1585), .D1(n1586), .SD(\adrram[2] ), .Z(n1592));
    L6MUX21 i1924 (.D0(n2021), .D1(n2022), .SD(\adrram[2] ), .Z(n2027));
    L6MUX21 i1736 (.D0(n1831), .D1(n1832), .SD(\adrram[2] ), .Z(n1839));
    L6MUX21 i1925 (.D0(n2023), .D1(n2024), .SD(\adrram[2] ), .Z(n2028));
    L6MUX21 i1737 (.D0(n1833), .D1(n1834), .SD(\adrram[2] ), .Z(n1840));
    L6MUX21 i1738 (.D0(n1835), .D1(n1836), .SD(\adrram[2] ), .Z(n1841));
    LUT4 i1464_3_lut (.A(\mem[0] [1]), .B(\mem[1] [1]), .C(\adrram[0] ), 
         .Z(n1567)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1464_3_lut.init = 16'hcaca;
    FD1P3AX mem_21__i0_i1 (.D(data[1]), .SP(we_N_63_enable_407), .CK(we_N_63), 
            .Q(\mem[21] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_21__i0_i1.GSR = "ENABLED";
    L6MUX21 i1550 (.D0(n1645), .D1(n1646), .SD(\adrram[2] ), .Z(n1653));
    L6MUX21 i1739 (.D0(n1837), .D1(n1838), .SD(\adrram[2] ), .Z(n1842));
    L6MUX21 i1551 (.D0(n1647), .D1(n1648), .SD(\adrram[2] ), .Z(n1654));
    L6MUX21 i1490 (.D0(n1587), .D1(n1588), .SD(\adrram[2] ), .Z(n1593));
    L6MUX21 i1552 (.D0(n1649), .D1(n1650), .SD(\adrram[2] ), .Z(n1655));
    L6MUX21 i1491 (.D0(n1589), .D1(n1590), .SD(\adrram[2] ), .Z(n1594));
    L6MUX21 i1553 (.D0(n1651), .D1(n1652), .SD(\adrram[2] ), .Z(n1656));
    L6MUX21 i1767 (.D0(n1862), .D1(n1863), .SD(\adrram[2] ), .Z(n1870));
    LUT4 i1748_3_lut (.A(\mem[42] [5]), .B(\mem[43] [5]), .C(\adrram[0] ), 
         .Z(n1851)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1748_3_lut.init = 16'hcaca;
    FD1P3AX mem_22__i0_i7 (.D(data[7]), .SP(we_N_63_enable_414), .CK(we_N_63), 
            .Q(\mem[22] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_22__i0_i7.GSR = "ENABLED";
    L6MUX21 i1860 (.D0(n1955), .D1(n1956), .SD(\adrram[2] ), .Z(n1963));
    PFUMX i1579 (.BLUT(n1672), .ALUT(n1673), .C0(\adrram[1] ), .Z(n1682));
    L6MUX21 i1768 (.D0(n1864), .D1(n1865), .SD(\adrram[2] ), .Z(n1871));
    L6MUX21 i1769 (.D0(n1866), .D1(n1867), .SD(\adrram[2] ), .Z(n1872));
    L6MUX21 i1861 (.D0(n1957), .D1(n1958), .SD(\adrram[2] ), .Z(n1964));
    L6MUX21 i1770 (.D0(n1868), .D1(n1869), .SD(\adrram[2] ), .Z(n1873));
    L6MUX21 i1862 (.D0(n1959), .D1(n1960), .SD(\adrram[2] ), .Z(n1965));
    L6MUX21 i1863 (.D0(n1961), .D1(n1962), .SD(\adrram[2] ), .Z(n1966));
    LUT4 i1747_3_lut (.A(\mem[40] [5]), .B(\mem[41] [5]), .C(\adrram[0] ), 
         .Z(n1850)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1747_3_lut.init = 16'hcaca;
    FD1P3AX mem_22__i0_i6 (.D(data[6]), .SP(we_N_63_enable_414), .CK(we_N_63), 
            .Q(\mem[22] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_22__i0_i6.GSR = "ENABLED";
    L6MUX21 i1612 (.D0(n1707), .D1(n1708), .SD(\adrram[2] ), .Z(n1715));
    L6MUX21 i1613 (.D0(n1709), .D1(n1710), .SD(\adrram[2] ), .Z(n1716));
    L6MUX21 i1614 (.D0(n1711), .D1(n1712), .SD(\adrram[2] ), .Z(n1717));
    L6MUX21 i1615 (.D0(n1713), .D1(n1714), .SD(\adrram[2] ), .Z(n1718));
    L6MUX21 i1643 (.D0(n1738), .D1(n1739), .SD(\adrram[2] ), .Z(n1746));
    L6MUX21 i1644 (.D0(n1740), .D1(n1741), .SD(\adrram[2] ), .Z(n1747));
    LUT4 i1746_3_lut (.A(\mem[38] [5]), .B(\mem[39] [5]), .C(\adrram[0] ), 
         .Z(n1849)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1746_3_lut.init = 16'hcaca;
    FD1P3AX mem_22__i0_i5 (.D(data[5]), .SP(we_N_63_enable_414), .CK(we_N_63), 
            .Q(\mem[22] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_22__i0_i5.GSR = "ENABLED";
    L6MUX21 i1645 (.D0(n1742), .D1(n1743), .SD(\adrram[2] ), .Z(n1748));
    L6MUX21 i1798 (.D0(n1893), .D1(n1894), .SD(\adrram[2] ), .Z(n1901));
    L6MUX21 i1646 (.D0(n1744), .D1(n1745), .SD(\adrram[2] ), .Z(n1749));
    LUT4 i1745_3_lut (.A(\mem[36] [5]), .B(\mem[37] [5]), .C(\adrram[0] ), 
         .Z(n1848)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1745_3_lut.init = 16'hcaca;
    L6MUX21 i1799 (.D0(n1895), .D1(n1896), .SD(\adrram[2] ), .Z(n1902));
    L6MUX21 i1800 (.D0(n1897), .D1(n1898), .SD(\adrram[2] ), .Z(n1903));
    LUT4 i1845_3_lut (.A(\mem[50] [2]), .B(\mem[51] [2]), .C(\adrram[0] ), 
         .Z(n1948)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1845_3_lut.init = 16'hcaca;
    FD1P3AX mem_22__i0_i4 (.D(data[4]), .SP(we_N_63_enable_414), .CK(we_N_63), 
            .Q(\mem[22] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_22__i0_i4.GSR = "ENABLED";
    L6MUX21 i1801 (.D0(n1899), .D1(n1900), .SD(\adrram[2] ), .Z(n1904));
    L6MUX21 i1674 (.D0(n1769), .D1(n1770), .SD(\adrram[2] ), .Z(n1777));
    L6MUX21 i1675 (.D0(n1771), .D1(n1772), .SD(\adrram[2] ), .Z(n1778));
    L6MUX21 i1676 (.D0(n1773), .D1(n1774), .SD(\adrram[2] ), .Z(n1779));
    LUT4 i1844_3_lut (.A(\mem[48] [2]), .B(\mem[49] [2]), .C(\adrram[0] ), 
         .Z(n1947)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1844_3_lut.init = 16'hcaca;
    L6MUX21 i1677 (.D0(n1775), .D1(n1776), .SD(\adrram[2] ), .Z(n1780));
    PFUMX i1511 (.BLUT(n1598), .ALUT(n1599), .C0(\adrram[1] ), .Z(n1614));
    LUT4 i1744_3_lut (.A(\mem[34] [5]), .B(\mem[35] [5]), .C(\adrram[0] ), 
         .Z(n1847)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1744_3_lut.init = 16'hcaca;
    FD1P3AX mem_22__i0_i3 (.D(data[3]), .SP(we_N_63_enable_414), .CK(we_N_63), 
            .Q(\mem[22] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_22__i0_i3.GSR = "ENABLED";
    PFUMX i1512 (.BLUT(n1600), .ALUT(n1601), .C0(\adrram[1] ), .Z(n1615));
    PFUMX i1513 (.BLUT(n1602), .ALUT(n1603), .C0(\adrram[1] ), .Z(n1616));
    LUT4 i1743_3_lut (.A(\mem[32] [5]), .B(\mem[33] [5]), .C(\adrram[0] ), 
         .Z(n1846)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1743_3_lut.init = 16'hcaca;
    FD1P3AX mem_22__i0_i2 (.D(data[2]), .SP(we_N_63_enable_414), .CK(we_N_63), 
            .Q(\mem[22] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_22__i0_i2.GSR = "ENABLED";
    PFUMX i1514 (.BLUT(n1604), .ALUT(n1605), .C0(\adrram[1] ), .Z(n1617));
    PFUMX i1454 (.BLUT(n1546), .ALUT(n1547), .C0(\adrram[1] ), .Z(n1557));
    LUT4 i1843_3_lut (.A(\mem[46] [2]), .B(\mem[47] [2]), .C(\adrram[0] ), 
         .Z(n1946)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1843_3_lut.init = 16'hcaca;
    FD1P3AX mem_22__i0_i1 (.D(data[1]), .SP(we_N_63_enable_414), .CK(we_N_63), 
            .Q(\mem[22] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_22__i0_i1.GSR = "ENABLED";
    PFUMX i1919 (.BLUT(n2011), .ALUT(n2012), .C0(\adrram[1] ), .Z(n2022));
    PFUMX i1886 (.BLUT(n1976), .ALUT(n1977), .C0(\adrram[1] ), .Z(n1989));
    LUT4 i1842_3_lut (.A(\mem[44] [2]), .B(\mem[45] [2]), .C(\adrram[0] ), 
         .Z(n1945)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1842_3_lut.init = 16'hcaca;
    FD1P3AX mem_47__i0_i2 (.D(data[2]), .SP(we_N_63_enable_416), .CK(we_N_63), 
            .Q(\mem[47] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_47__i0_i2.GSR = "ENABLED";
    PFUMX i1515 (.BLUT(n1606), .ALUT(n1607), .C0(\adrram[1] ), .Z(n1618));
    PFUMX i1516 (.BLUT(n1608), .ALUT(n1609), .C0(\adrram[1] ), .Z(n1619));
    LUT4 i1841_3_lut (.A(\mem[42] [2]), .B(\mem[43] [2]), .C(\adrram[0] ), 
         .Z(n1944)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1841_3_lut.init = 16'hcaca;
    LUT4 i1840_3_lut (.A(\mem[40] [2]), .B(\mem[41] [2]), .C(\adrram[0] ), 
         .Z(n1943)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1840_3_lut.init = 16'hcaca;
    PFUMX i1517 (.BLUT(n1610), .ALUT(n1611), .C0(\adrram[1] ), .Z(n1620));
    PFUMX i1518 (.BLUT(n1612), .ALUT(n1613), .C0(\adrram[1] ), .Z(n1621));
    LUT4 i1442_3_lut (.A(\mem[18] [0]), .B(\mem[19] [0]), .C(\adrram[0] ), 
         .Z(n1545)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1442_3_lut.init = 16'hcaca;
    LUT4 i1441_3_lut (.A(\mem[16] [0]), .B(\mem[17] [0]), .C(\adrram[0] ), 
         .Z(n1544)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1441_3_lut.init = 16'hcaca;
    PFUMX i1821 (.BLUT(n1908), .ALUT(n1909), .C0(\adrram[1] ), .Z(n1924));
    PFUMX i1887 (.BLUT(n1978), .ALUT(n1979), .C0(\adrram[1] ), .Z(n1990));
    LUT4 i1839_3_lut (.A(\mem[38] [2]), .B(\mem[39] [2]), .C(\adrram[0] ), 
         .Z(n1942)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1839_3_lut.init = 16'hcaca;
    LUT4 i1838_3_lut (.A(\mem[36] [2]), .B(\mem[37] [2]), .C(\adrram[0] ), 
         .Z(n1941)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1838_3_lut.init = 16'hcaca;
    PFUMX i1822 (.BLUT(n1910), .ALUT(n1911), .C0(\adrram[1] ), .Z(n1925));
    LUT4 i1837_3_lut (.A(\mem[34] [2]), .B(\mem[35] [2]), .C(\adrram[0] ), 
         .Z(n1940)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1837_3_lut.init = 16'hcaca;
    LUT4 i1836_3_lut (.A(\mem[32] [2]), .B(\mem[33] [2]), .C(\adrram[0] ), 
         .Z(n1939)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1836_3_lut.init = 16'hcaca;
    LUT4 i1440_3_lut (.A(\mem[14] [0]), .B(\mem[15] [0]), .C(\adrram[0] ), 
         .Z(n1543)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1440_3_lut.init = 16'hcaca;
    LUT4 i1439_3_lut (.A(\mem[12] [0]), .B(\mem[13] [0]), .C(\adrram[0] ), 
         .Z(n1542)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1439_3_lut.init = 16'hcaca;
    LUT4 i1438_3_lut (.A(\mem[10] [0]), .B(\mem[11] [0]), .C(\adrram[0] ), 
         .Z(n1541)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1438_3_lut.init = 16'hcaca;
    LUT4 i1437_3_lut (.A(\mem[8] [0]), .B(\mem[9] [0]), .C(\adrram[0] ), 
         .Z(n1540)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1437_3_lut.init = 16'hcaca;
    PFUMX i1823 (.BLUT(n1912), .ALUT(n1913), .C0(\adrram[1] ), .Z(n1926));
    PFUMX i1920 (.BLUT(n2013), .ALUT(n2014), .C0(\adrram[1] ), .Z(n2023));
    LUT4 i1541_3_lut (.A(\mem[30] [3]), .B(\mem[31] [3]), .C(\adrram[0] ), 
         .Z(n1644)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1541_3_lut.init = 16'hcaca;
    FD1P3AX mem_47__i0_i1 (.D(data[1]), .SP(we_N_63_enable_416), .CK(we_N_63), 
            .Q(\mem[47] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_47__i0_i1.GSR = "ENABLED";
    PFUMX i1888 (.BLUT(n1980), .ALUT(n1981), .C0(\adrram[1] ), .Z(n1991));
    LUT4 i1540_3_lut (.A(\mem[28] [3]), .B(\mem[29] [3]), .C(\adrram[0] ), 
         .Z(n1643)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1540_3_lut.init = 16'hcaca;
    PFUMX i1824 (.BLUT(n1914), .ALUT(n1915), .C0(\adrram[1] ), .Z(n1927));
    LUT4 i1539_3_lut (.A(\mem[26] [3]), .B(\mem[27] [3]), .C(\adrram[0] ), 
         .Z(n1642)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1539_3_lut.init = 16'hcaca;
    LUT4 i1538_3_lut (.A(\mem[24] [3]), .B(\mem[25] [3]), .C(\adrram[0] ), 
         .Z(n1641)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1538_3_lut.init = 16'hcaca;
    FD1P3AX mem_46__i0_i7 (.D(data[7]), .SP(we_N_63_enable_423), .CK(we_N_63), 
            .Q(\mem[46] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_46__i0_i7.GSR = "ENABLED";
    PFUMX i1697 (.BLUT(n1784), .ALUT(n1785), .C0(\adrram[1] ), .Z(n1800));
    LUT4 i1537_3_lut (.A(\mem[22] [3]), .B(\mem[23] [3]), .C(\adrram[0] ), 
         .Z(n1640)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1537_3_lut.init = 16'hcaca;
    LUT4 i1536_3_lut (.A(\mem[20] [3]), .B(\mem[21] [3]), .C(\adrram[0] ), 
         .Z(n1639)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1536_3_lut.init = 16'hcaca;
    PFUMX i1825 (.BLUT(n1916), .ALUT(n1917), .C0(\adrram[1] ), .Z(n1928));
    LUT4 i1535_3_lut (.A(\mem[18] [3]), .B(\mem[19] [3]), .C(\adrram[0] ), 
         .Z(n1638)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1535_3_lut.init = 16'hcaca;
    FD1P3AX mem_46__i0_i6 (.D(data[6]), .SP(we_N_63_enable_423), .CK(we_N_63), 
            .Q(\mem[46] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_46__i0_i6.GSR = "ENABLED";
    PFUMX i1698 (.BLUT(n1786), .ALUT(n1787), .C0(\adrram[1] ), .Z(n1801));
    LUT4 i1534_3_lut (.A(\mem[16] [3]), .B(\mem[17] [3]), .C(\adrram[0] ), 
         .Z(n1637)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1534_3_lut.init = 16'hcaca;
    LUT4 i1533_3_lut (.A(\mem[14] [3]), .B(\mem[15] [3]), .C(\adrram[0] ), 
         .Z(n1636)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1533_3_lut.init = 16'hcaca;
    PFUMX i1699 (.BLUT(n1788), .ALUT(n1789), .C0(\adrram[1] ), .Z(n1802));
    PFUMX i1889 (.BLUT(n1982), .ALUT(n1983), .C0(\adrram[1] ), .Z(n1992));
    LUT4 i1532_3_lut (.A(\mem[12] [3]), .B(\mem[13] [3]), .C(\adrram[0] ), 
         .Z(n1635)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1532_3_lut.init = 16'hcaca;
    FD1P3AX mem_46__i0_i5 (.D(data[5]), .SP(we_N_63_enable_423), .CK(we_N_63), 
            .Q(\mem[46] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_46__i0_i5.GSR = "ENABLED";
    PFUMX i1486 (.BLUT(n1579), .ALUT(n1580), .C0(\adrram[1] ), .Z(n1589));
    LUT4 i1531_3_lut (.A(\mem[10] [3]), .B(\mem[11] [3]), .C(\adrram[0] ), 
         .Z(n1634)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1531_3_lut.init = 16'hcaca;
    PFUMX i1487 (.BLUT(n1581), .ALUT(n1582), .C0(\adrram[1] ), .Z(n1590));
    LUT4 i1530_3_lut (.A(\mem[8] [3]), .B(\mem[9] [3]), .C(\adrram[0] ), 
         .Z(n1633)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1530_3_lut.init = 16'hcaca;
    FD1P3AX mem_46__i0_i4 (.D(data[4]), .SP(we_N_63_enable_423), .CK(we_N_63), 
            .Q(\mem[46] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_46__i0_i4.GSR = "ENABLED";
    LUT4 i1727_3_lut (.A(\mem[62] [6]), .B(\mem[63] [6]), .C(\adrram[0] ), 
         .Z(n1830)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1727_3_lut.init = 16'hcaca;
    PFUMX i1728 (.BLUT(n1815), .ALUT(n1816), .C0(\adrram[1] ), .Z(n1831));
    LUT4 i1726_3_lut (.A(\mem[60] [6]), .B(\mem[61] [6]), .C(\adrram[0] ), 
         .Z(n1829)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1726_3_lut.init = 16'hcaca;
    PFUMX i1729 (.BLUT(n1817), .ALUT(n1818), .C0(\adrram[1] ), .Z(n1832));
    PFUMX i1730 (.BLUT(n1819), .ALUT(n1820), .C0(\adrram[1] ), .Z(n1833));
    LUT4 i1529_3_lut (.A(\mem[6] [3]), .B(\mem[7] [3]), .C(\adrram[0] ), 
         .Z(n1632)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1529_3_lut.init = 16'hcaca;
    FD1P3AX mem_46__i0_i3 (.D(data[3]), .SP(we_N_63_enable_423), .CK(we_N_63), 
            .Q(\mem[46] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_46__i0_i3.GSR = "ENABLED";
    LUT4 i1528_3_lut (.A(\mem[4] [3]), .B(\mem[5] [3]), .C(\adrram[0] ), 
         .Z(n1631)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1528_3_lut.init = 16'hcaca;
    PFUMX i1857 (.BLUT(n1949), .ALUT(n1950), .C0(\adrram[1] ), .Z(n1960));
    LUT4 i1436_3_lut (.A(\mem[6] [0]), .B(\mem[7] [0]), .C(\adrram[0] ), 
         .Z(n1539)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1436_3_lut.init = 16'hcaca;
    LUT4 i1905_3_lut (.A(\mem[46] [0]), .B(\mem[47] [0]), .C(\adrram[0] ), 
         .Z(n2008)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1905_3_lut.init = 16'hcaca;
    PFUMX i1483 (.BLUT(n1573), .ALUT(n1574), .C0(\adrram[1] ), .Z(n1586));
    LUT4 i1435_3_lut (.A(\mem[4] [0]), .B(\mem[5] [0]), .C(\adrram[0] ), 
         .Z(n1538)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1435_3_lut.init = 16'hcaca;
    FD1P3AX mem_46__i0_i2 (.D(data[2]), .SP(we_N_63_enable_423), .CK(we_N_63), 
            .Q(\mem[46] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_46__i0_i2.GSR = "ENABLED";
    LUT4 i1627_3_lut (.A(\mem[16] [6]), .B(\mem[17] [6]), .C(\adrram[0] ), 
         .Z(n1730)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1627_3_lut.init = 16'hcaca;
    PFUMX i1762 (.BLUT(n1852), .ALUT(n1853), .C0(\adrram[1] ), .Z(n1865));
    LUT4 i1904_3_lut (.A(\mem[44] [0]), .B(\mem[45] [0]), .C(\adrram[0] ), 
         .Z(n2007)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1904_3_lut.init = 16'hcaca;
    PFUMX i1573 (.BLUT(n1660), .ALUT(n1661), .C0(\adrram[1] ), .Z(n1676));
    LUT4 i1901_3_lut (.A(\mem[38] [0]), .B(\mem[39] [0]), .C(\adrram[0] ), 
         .Z(n2004)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1901_3_lut.init = 16'hcaca;
    FD1P3AX mem_46__i0_i1 (.D(data[1]), .SP(we_N_63_enable_423), .CK(we_N_63), 
            .Q(\mem[46] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_46__i0_i1.GSR = "ENABLED";
    LUT4 i1626_3_lut (.A(\mem[14] [6]), .B(\mem[15] [6]), .C(\adrram[0] ), 
         .Z(n1729)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1626_3_lut.init = 16'hcaca;
    PFUMX i1481 (.BLUT(n1569), .ALUT(n1570), .C0(\adrram[1] ), .Z(n1584));
    LUT4 i1868_3_lut (.A(\mem[34] [1]), .B(\mem[35] [1]), .C(\adrram[0] ), 
         .Z(n1971)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1868_3_lut.init = 16'hcaca;
    PFUMX i1858 (.BLUT(n1951), .ALUT(n1952), .C0(\adrram[1] ), .Z(n1961));
    LUT4 i1900_3_lut (.A(\mem[36] [0]), .B(\mem[37] [0]), .C(\adrram[0] ), 
         .Z(n2003)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1900_3_lut.init = 16'hcaca;
    PFUMX i1482 (.BLUT(n1571), .ALUT(n1572), .C0(\adrram[1] ), .Z(n1585));
    LUT4 i1625_3_lut (.A(\mem[12] [6]), .B(\mem[13] [6]), .C(\adrram[0] ), 
         .Z(n1728)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1625_3_lut.init = 16'hcaca;
    PFUMX i1764 (.BLUT(n1856), .ALUT(n1857), .C0(\adrram[1] ), .Z(n1867));
    LUT4 i1777_3_lut (.A(\mem[38] [4]), .B(\mem[39] [4]), .C(\adrram[0] ), 
         .Z(n1880)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1777_3_lut.init = 16'hcaca;
    LUT4 i1595_3_lut (.A(\mem[14] [5]), .B(\mem[15] [5]), .C(\adrram[0] ), 
         .Z(n1698)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1595_3_lut.init = 16'hcaca;
    LUT4 i2222_2_lut_2_lut_3_lut_4_lut (.A(\adrram[1] ), .B(n2250), .C(n2249), 
         .D(\adrram[3] ), .Z(we_N_63_enable_322)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2222_2_lut_2_lut_3_lut_4_lut.init = 16'h0200;
    PFUMX i1731 (.BLUT(n1821), .ALUT(n1822), .C0(\adrram[1] ), .Z(n1834));
    LUT4 i1867_3_lut (.A(\mem[32] [1]), .B(\mem[33] [1]), .C(\adrram[0] ), 
         .Z(n1970)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1867_3_lut.init = 16'hcaca;
    LUT4 i1776_3_lut (.A(\mem[36] [4]), .B(\mem[37] [4]), .C(\adrram[0] ), 
         .Z(n1879)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1776_3_lut.init = 16'hcaca;
    LUT4 i1434_3_lut (.A(\mem[2] [0]), .B(\mem[3] [0]), .C(\adrram[0] ), 
         .Z(n1537)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1434_3_lut.init = 16'hcaca;
    FD1P3AX mem_45__i0_i7 (.D(data[7]), .SP(we_N_63_enable_446), .CK(we_N_63), 
            .Q(\mem[45] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_45__i0_i7.GSR = "ENABLED";
    LUT4 i1783_3_lut (.A(\mem[50] [4]), .B(\mem[51] [4]), .C(\adrram[0] ), 
         .Z(n1886)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1783_3_lut.init = 16'hcaca;
    FD1P3AX mem_45__i0_i6 (.D(data[6]), .SP(we_N_63_enable_446), .CK(we_N_63), 
            .Q(\mem[45] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_45__i0_i6.GSR = "ENABLED";
    LUT4 i1594_3_lut (.A(\mem[12] [5]), .B(\mem[13] [5]), .C(\adrram[0] ), 
         .Z(n1697)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1594_3_lut.init = 16'hcaca;
    FD1P3AY mem_62__i0_i7 (.D(data[7]), .SP(we_N_63_enable_433), .CK(we_N_63), 
            .Q(\mem[62] [7])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_62__i0_i7.GSR = "ENABLED";
    FD1P3AY mem_62__i0_i6 (.D(data[6]), .SP(we_N_63_enable_433), .CK(we_N_63), 
            .Q(\mem[62] [6])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_62__i0_i6.GSR = "ENABLED";
    FD1P3AY mem_62__i0_i5 (.D(data[5]), .SP(we_N_63_enable_433), .CK(we_N_63), 
            .Q(\mem[62] [5])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_62__i0_i5.GSR = "ENABLED";
    FD1P3AY mem_62__i0_i4 (.D(data[4]), .SP(we_N_63_enable_433), .CK(we_N_63), 
            .Q(\mem[62] [4])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_62__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_45__i0_i5 (.D(data[5]), .SP(we_N_63_enable_446), .CK(we_N_63), 
            .Q(\mem[45] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_45__i0_i5.GSR = "ENABLED";
    LUT4 i1563_3_lut (.A(\mem[12] [4]), .B(\mem[13] [4]), .C(\adrram[0] ), 
         .Z(n1666)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1563_3_lut.init = 16'hcaca;
    FD1P3AY mem_62__i0_i3 (.D(data[3]), .SP(we_N_63_enable_433), .CK(we_N_63), 
            .Q(\mem[62] [3])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_62__i0_i3.GSR = "ENABLED";
    FD1P3AY mem_62__i0_i2 (.D(data[2]), .SP(we_N_63_enable_433), .CK(we_N_63), 
            .Q(\mem[62] [2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_62__i0_i2.GSR = "ENABLED";
    FD1P3AY mem_62__i0_i1 (.D(data[1]), .SP(we_N_63_enable_433), .CK(we_N_63), 
            .Q(\mem[62] [1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_62__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_61__i0_i7 (.D(data[7]), .SP(we_N_63_enable_443), .CK(we_N_63), 
            .Q(\mem[61] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_61__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_45__i0_i4 (.D(data[4]), .SP(we_N_63_enable_446), .CK(we_N_63), 
            .Q(\mem[45] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_45__i0_i4.GSR = "ENABLED";
    LUT4 i1665_3_lut (.A(\mem[30] [7]), .B(\mem[31] [7]), .C(\adrram[0] ), 
         .Z(n1768)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1665_3_lut.init = 16'hcaca;
    FD1P3AX mem_61__i0_i6 (.D(data[6]), .SP(we_N_63_enable_443), .CK(we_N_63), 
            .Q(\mem[61] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_61__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_61__i0_i5 (.D(data[5]), .SP(we_N_63_enable_443), .CK(we_N_63), 
            .Q(\mem[61] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_61__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_61__i0_i4 (.D(data[4]), .SP(we_N_63_enable_443), .CK(we_N_63), 
            .Q(\mem[61] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_61__i0_i4.GSR = "ENABLED";
    LUT4 i1433_3_lut (.A(\mem[0] [0]), .B(\mem[1] [0]), .C(\adrram[0] ), 
         .Z(n1536)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1433_3_lut.init = 16'hcaca;
    FD1P3AX mem_45__i0_i3 (.D(data[3]), .SP(we_N_63_enable_446), .CK(we_N_63), 
            .Q(\mem[45] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_45__i0_i3.GSR = "ENABLED";
    LUT4 i1782_3_lut (.A(\mem[48] [4]), .B(\mem[49] [4]), .C(\adrram[0] ), 
         .Z(n1885)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1782_3_lut.init = 16'hcaca;
    LUT4 i1775_3_lut (.A(\mem[34] [4]), .B(\mem[35] [4]), .C(\adrram[0] ), 
         .Z(n1878)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1775_3_lut.init = 16'hcaca;
    FD1P3AX mem_61__i0_i3 (.D(data[3]), .SP(we_N_63_enable_443), .CK(we_N_63), 
            .Q(\mem[61] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_61__i0_i3.GSR = "ENABLED";
    LUT4 i1664_3_lut (.A(\mem[28] [7]), .B(\mem[29] [7]), .C(\adrram[0] ), 
         .Z(n1767)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1664_3_lut.init = 16'hcaca;
    FD1P3AX mem_61__i0_i2 (.D(data[2]), .SP(we_N_63_enable_443), .CK(we_N_63), 
            .Q(\mem[61] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_61__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_45__i0_i2 (.D(data[2]), .SP(we_N_63_enable_446), .CK(we_N_63), 
            .Q(\mem[45] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_45__i0_i2.GSR = "ENABLED";
    LUT4 i1774_3_lut (.A(\mem[32] [4]), .B(\mem[33] [4]), .C(\adrram[0] ), 
         .Z(n1877)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1774_3_lut.init = 16'hcaca;
    FD1P3AX mem_61__i0_i1 (.D(data[1]), .SP(we_N_63_enable_443), .CK(we_N_63), 
            .Q(\mem[61] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_61__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_60__i0_i7 (.D(data[7]), .SP(we_N_63_enable_452), .CK(we_N_63), 
            .Q(\mem[60] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_60__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_60__i0_i6 (.D(data[6]), .SP(we_N_63_enable_452), .CK(we_N_63), 
            .Q(\mem[60] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_60__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_45__i0_i1 (.D(data[1]), .SP(we_N_63_enable_446), .CK(we_N_63), 
            .Q(\mem[45] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_45__i0_i1.GSR = "ENABLED";
    LUT4 i1593_3_lut (.A(\mem[10] [5]), .B(\mem[11] [5]), .C(\adrram[0] ), 
         .Z(n1696)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1593_3_lut.init = 16'hcaca;
    FD1P3AX mem_60__i0_i5 (.D(data[5]), .SP(we_N_63_enable_452), .CK(we_N_63), 
            .Q(\mem[60] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_60__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_60__i0_i4 (.D(data[4]), .SP(we_N_63_enable_452), .CK(we_N_63), 
            .Q(\mem[60] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_60__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_60__i0_i3 (.D(data[3]), .SP(we_N_63_enable_452), .CK(we_N_63), 
            .Q(\mem[60] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_60__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_44__i0_i7 (.D(data[7]), .SP(we_N_63_enable_475), .CK(we_N_63), 
            .Q(\mem[44] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_44__i0_i7.GSR = "ENABLED";
    LUT4 i1757_3_lut (.A(\mem[60] [5]), .B(\mem[61] [5]), .C(\adrram[0] ), 
         .Z(n1860)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1757_3_lut.init = 16'hcaca;
    FD1P3AX mem_60__i0_i2 (.D(data[2]), .SP(we_N_63_enable_452), .CK(we_N_63), 
            .Q(\mem[60] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_60__i0_i2.GSR = "ENABLED";
    LUT4 i1448_3_lut (.A(\mem[30] [0]), .B(\mem[31] [0]), .C(\adrram[0] ), 
         .Z(n1551)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1448_3_lut.init = 16'hcaca;
    FD1P3AX mem_60__i0_i1 (.D(data[1]), .SP(we_N_63_enable_452), .CK(we_N_63), 
            .Q(\mem[60] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_60__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_44__i0_i6 (.D(data[6]), .SP(we_N_63_enable_475), .CK(we_N_63), 
            .Q(\mem[44] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_44__i0_i6.GSR = "ENABLED";
    LUT4 i1624_3_lut (.A(\mem[10] [6]), .B(\mem[11] [6]), .C(\adrram[0] ), 
         .Z(n1727)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1624_3_lut.init = 16'hcaca;
    LUT4 i1592_3_lut (.A(\mem[8] [5]), .B(\mem[9] [5]), .C(\adrram[0] ), 
         .Z(n1695)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1592_3_lut.init = 16'hcaca;
    LUT4 i1562_3_lut (.A(\mem[10] [4]), .B(\mem[11] [4]), .C(\adrram[0] ), 
         .Z(n1665)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1562_3_lut.init = 16'hcaca;
    LUT4 i1752_3_lut (.A(\mem[50] [5]), .B(\mem[51] [5]), .C(\adrram[0] ), 
         .Z(n1855)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1752_3_lut.init = 16'hcaca;
    LUT4 i2191_2_lut_2_lut_3_lut_4_lut (.A(\adrram[1] ), .B(n2250), .C(n2248), 
         .D(\adrram[3] ), .Z(we_N_63_enable_175)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2191_2_lut_2_lut_3_lut_4_lut.init = 16'h0002;
    LUT4 i1663_3_lut (.A(\mem[26] [7]), .B(\mem[27] [7]), .C(\adrram[0] ), 
         .Z(n1766)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1663_3_lut.init = 16'hcaca;
    FD1P3AX mem_59__i0_i7 (.D(data[7]), .SP(we_N_63_enable_461), .CK(we_N_63), 
            .Q(\mem[59] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_59__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_59__i0_i6 (.D(data[6]), .SP(we_N_63_enable_461), .CK(we_N_63), 
            .Q(\mem[59] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_59__i0_i6.GSR = "ENABLED";
    LUT4 i1447_3_lut (.A(\mem[28] [0]), .B(\mem[29] [0]), .C(\adrram[0] ), 
         .Z(n1550)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1447_3_lut.init = 16'hcaca;
    FD1P3AX mem_59__i0_i5 (.D(data[5]), .SP(we_N_63_enable_461), .CK(we_N_63), 
            .Q(\mem[59] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_59__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_44__i0_i5 (.D(data[5]), .SP(we_N_63_enable_475), .CK(we_N_63), 
            .Q(\mem[44] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_44__i0_i5.GSR = "ENABLED";
    LUT4 i1623_3_lut (.A(\mem[8] [6]), .B(\mem[9] [6]), .C(\adrram[0] ), 
         .Z(n1726)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1623_3_lut.init = 16'hcaca;
    LUT4 i1603_3_lut (.A(\mem[30] [5]), .B(\mem[31] [5]), .C(\adrram[0] ), 
         .Z(n1706)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1603_3_lut.init = 16'hcaca;
    LUT4 i1561_3_lut (.A(\mem[8] [4]), .B(\mem[9] [4]), .C(\adrram[0] ), 
         .Z(n1664)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1561_3_lut.init = 16'hcaca;
    LUT4 i1851_3_lut (.A(\mem[62] [2]), .B(\mem[63] [2]), .C(\adrram[0] ), 
         .Z(n1954)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1851_3_lut.init = 16'hcaca;
    LUT4 i1662_3_lut (.A(\mem[24] [7]), .B(\mem[25] [7]), .C(\adrram[0] ), 
         .Z(n1765)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1662_3_lut.init = 16'hcaca;
    LUT4 i1602_3_lut (.A(\mem[28] [5]), .B(\mem[29] [5]), .C(\adrram[0] ), 
         .Z(n1705)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1602_3_lut.init = 16'hcaca;
    FD1P3AX mem_59__i0_i4 (.D(data[4]), .SP(we_N_63_enable_461), .CK(we_N_63), 
            .Q(\mem[59] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_59__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_59__i0_i3 (.D(data[3]), .SP(we_N_63_enable_461), .CK(we_N_63), 
            .Q(\mem[59] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_59__i0_i3.GSR = "ENABLED";
    LUT4 i1591_3_lut (.A(\mem[6] [5]), .B(\mem[7] [5]), .C(\adrram[0] ), 
         .Z(n1694)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1591_3_lut.init = 16'hcaca;
    FD1P3AX mem_59__i0_i2 (.D(data[2]), .SP(we_N_63_enable_461), .CK(we_N_63), 
            .Q(\mem[59] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_59__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_59__i0_i1 (.D(data[1]), .SP(we_N_63_enable_461), .CK(we_N_63), 
            .Q(\mem[59] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_59__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_44__i0_i4 (.D(data[4]), .SP(we_N_63_enable_475), .CK(we_N_63), 
            .Q(\mem[44] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_44__i0_i4.GSR = "ENABLED";
    LUT4 i1850_3_lut (.A(\mem[60] [2]), .B(\mem[61] [2]), .C(\adrram[0] ), 
         .Z(n1953)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1850_3_lut.init = 16'hcaca;
    LUT4 i1751_3_lut (.A(\mem[48] [5]), .B(\mem[49] [5]), .C(\adrram[0] ), 
         .Z(n1854)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1751_3_lut.init = 16'hcaca;
    LUT4 i1899_3_lut (.A(\mem[34] [0]), .B(\mem[35] [0]), .C(\adrram[0] ), 
         .Z(n2002)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1899_3_lut.init = 16'hcaca;
    LUT4 i1661_3_lut (.A(\mem[22] [7]), .B(\mem[23] [7]), .C(\adrram[0] ), 
         .Z(n1764)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1661_3_lut.init = 16'hcaca;
    LUT4 i1898_3_lut (.A(\mem[32] [0]), .B(\mem[33] [0]), .C(\adrram[0] ), 
         .Z(n2001)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1898_3_lut.init = 16'hcaca;
    FD1P3AX mem_58__i0_i7 (.D(data[7]), .SP(we_N_63_enable_470), .CK(we_N_63), 
            .Q(\mem[58] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_58__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_58__i0_i6 (.D(data[6]), .SP(we_N_63_enable_470), .CK(we_N_63), 
            .Q(\mem[58] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_58__i0_i6.GSR = "ENABLED";
    LUT4 i1622_3_lut (.A(\mem[6] [6]), .B(\mem[7] [6]), .C(\adrram[0] ), 
         .Z(n1725)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1622_3_lut.init = 16'hcaca;
    FD1P3AX mem_58__i0_i5 (.D(data[5]), .SP(we_N_63_enable_470), .CK(we_N_63), 
            .Q(\mem[58] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_58__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_58__i0_i4 (.D(data[4]), .SP(we_N_63_enable_470), .CK(we_N_63), 
            .Q(\mem[58] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_58__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_44__i0_i3 (.D(data[3]), .SP(we_N_63_enable_475), .CK(we_N_63), 
            .Q(\mem[44] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_44__i0_i3.GSR = "ENABLED";
    LUT4 i1660_3_lut (.A(\mem[20] [7]), .B(\mem[21] [7]), .C(\adrram[0] ), 
         .Z(n1763)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1660_3_lut.init = 16'hcaca;
    FD1P3AX mem_58__i0_i3 (.D(data[3]), .SP(we_N_63_enable_470), .CK(we_N_63), 
            .Q(\mem[58] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_58__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_58__i0_i2 (.D(data[2]), .SP(we_N_63_enable_470), .CK(we_N_63), 
            .Q(\mem[58] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_58__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_58__i0_i1 (.D(data[1]), .SP(we_N_63_enable_470), .CK(we_N_63), 
            .Q(\mem[58] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_58__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_44__i0_i2 (.D(data[2]), .SP(we_N_63_enable_475), .CK(we_N_63), 
            .Q(\mem[44] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_44__i0_i2.GSR = "ENABLED";
    LUT4 i1789_3_lut (.A(\mem[62] [4]), .B(\mem[63] [4]), .C(\adrram[0] ), 
         .Z(n1892)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1789_3_lut.init = 16'hcaca;
    LUT4 i1621_3_lut (.A(\mem[4] [6]), .B(\mem[5] [6]), .C(\adrram[0] ), 
         .Z(n1724)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1621_3_lut.init = 16'hcaca;
    LUT4 i1788_3_lut (.A(\mem[60] [4]), .B(\mem[61] [4]), .C(\adrram[0] ), 
         .Z(n1891)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1788_3_lut.init = 16'hcaca;
    LUT4 i1659_3_lut (.A(\mem[18] [7]), .B(\mem[19] [7]), .C(\adrram[0] ), 
         .Z(n1762)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1659_3_lut.init = 16'hcaca;
    FD1P3AX mem_57__i0_i7 (.D(data[7]), .SP(we_N_63_enable_479), .CK(we_N_63), 
            .Q(\mem[57] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_57__i0_i7.GSR = "ENABLED";
    LUT4 i1658_3_lut (.A(\mem[16] [7]), .B(\mem[17] [7]), .C(\adrram[0] ), 
         .Z(n1761)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1658_3_lut.init = 16'hcaca;
    FD1P3AX mem_57__i0_i6 (.D(data[6]), .SP(we_N_63_enable_479), .CK(we_N_63), 
            .Q(\mem[57] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_57__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_57__i0_i5 (.D(data[5]), .SP(we_N_63_enable_479), .CK(we_N_63), 
            .Q(\mem[57] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_57__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_44__i0_i1 (.D(data[1]), .SP(we_N_63_enable_475), .CK(we_N_63), 
            .Q(\mem[44] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_44__i0_i1.GSR = "ENABLED";
    LUT4 i1634_3_lut (.A(\mem[30] [6]), .B(\mem[31] [6]), .C(\adrram[0] ), 
         .Z(n1737)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1634_3_lut.init = 16'hcaca;
    LUT4 i1657_3_lut (.A(\mem[14] [7]), .B(\mem[15] [7]), .C(\adrram[0] ), 
         .Z(n1760)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1657_3_lut.init = 16'hcaca;
    LUT4 i1633_3_lut (.A(\mem[28] [6]), .B(\mem[29] [6]), .C(\adrram[0] ), 
         .Z(n1736)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1633_3_lut.init = 16'hcaca;
    LUT4 i1781_3_lut (.A(\mem[46] [4]), .B(\mem[47] [4]), .C(\adrram[0] ), 
         .Z(n1884)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1781_3_lut.init = 16'hcaca;
    FD1P3AX mem_57__i0_i4 (.D(data[4]), .SP(we_N_63_enable_479), .CK(we_N_63), 
            .Q(\mem[57] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_57__i0_i4.GSR = "ENABLED";
    PFUMX i1732 (.BLUT(n1823), .ALUT(n1824), .C0(\adrram[1] ), .Z(n1835));
    FD1P3AX mem_57__i0_i3 (.D(data[3]), .SP(we_N_63_enable_479), .CK(we_N_63), 
            .Q(\mem[57] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_57__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_57__i0_i2 (.D(data[2]), .SP(we_N_63_enable_479), .CK(we_N_63), 
            .Q(\mem[57] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_57__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_57__i0_i1 (.D(data[1]), .SP(we_N_63_enable_479), .CK(we_N_63), 
            .Q(\mem[57] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_57__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_43__i0_i7 (.D(data[7]), .SP(we_N_63_enable_511), .CK(we_N_63), 
            .Q(\mem[43] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_43__i0_i7.GSR = "ENABLED";
    PFUMX i1733 (.BLUT(n1825), .ALUT(n1826), .C0(\adrram[1] ), .Z(n1836));
    LUT4 i1601_3_lut (.A(\mem[26] [5]), .B(\mem[27] [5]), .C(\adrram[0] ), 
         .Z(n1704)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1601_3_lut.init = 16'hcaca;
    FD1P3AX mem_56__i0_i7 (.D(data[7]), .SP(we_N_63_enable_488), .CK(we_N_63), 
            .Q(\mem[56] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_56__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_56__i0_i6 (.D(data[6]), .SP(we_N_63_enable_488), .CK(we_N_63), 
            .Q(\mem[56] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_56__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_56__i0_i5 (.D(data[5]), .SP(we_N_63_enable_488), .CK(we_N_63), 
            .Q(\mem[56] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_56__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_56__i0_i4 (.D(data[4]), .SP(we_N_63_enable_488), .CK(we_N_63), 
            .Q(\mem[56] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_56__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_43__i0_i6 (.D(data[6]), .SP(we_N_63_enable_511), .CK(we_N_63), 
            .Q(\mem[43] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_43__i0_i6.GSR = "ENABLED";
    PFUMX i1734 (.BLUT(n1827), .ALUT(n1828), .C0(\adrram[1] ), .Z(n1837));
    PFUMX i1542 (.BLUT(n1629), .ALUT(n1630), .C0(\adrram[1] ), .Z(n1645));
    LUT4 i1590_3_lut (.A(\mem[4] [5]), .B(\mem[5] [5]), .C(\adrram[0] ), 
         .Z(n1693)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1590_3_lut.init = 16'hcaca;
    FD1P3AX mem_56__i0_i3 (.D(data[3]), .SP(we_N_63_enable_488), .CK(we_N_63), 
            .Q(\mem[56] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_56__i0_i3.GSR = "ENABLED";
    PFUMX i1484 (.BLUT(n1575), .ALUT(n1576), .C0(\adrram[1] ), .Z(n1587));
    FD1P3AX mem_56__i0_i2 (.D(data[2]), .SP(we_N_63_enable_488), .CK(we_N_63), 
            .Q(\mem[56] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_56__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_56__i0_i1 (.D(data[1]), .SP(we_N_63_enable_488), .CK(we_N_63), 
            .Q(\mem[56] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_56__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_43__i0_i5 (.D(data[5]), .SP(we_N_63_enable_511), .CK(we_N_63), 
            .Q(\mem[43] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_43__i0_i5.GSR = "ENABLED";
    PFUMX i1765 (.BLUT(n1858), .ALUT(n1859), .C0(\adrram[1] ), .Z(n1868));
    FD1P3AX mem_55__i0_i7 (.D(data[7]), .SP(we_N_63_enable_497), .CK(we_N_63), 
            .Q(\mem[55] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_55__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_55__i0_i6 (.D(data[6]), .SP(we_N_63_enable_497), .CK(we_N_63), 
            .Q(\mem[55] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_55__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_55__i0_i5 (.D(data[5]), .SP(we_N_63_enable_497), .CK(we_N_63), 
            .Q(\mem[55] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_55__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_55__i0_i4 (.D(data[4]), .SP(we_N_63_enable_497), .CK(we_N_63), 
            .Q(\mem[55] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_55__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_43__i0_i4 (.D(data[4]), .SP(we_N_63_enable_511), .CK(we_N_63), 
            .Q(\mem[43] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_43__i0_i4.GSR = "ENABLED";
    PFUMX i1577 (.BLUT(n1668), .ALUT(n1669), .C0(\adrram[1] ), .Z(n1680));
    PFUMX i1608 (.BLUT(n1699), .ALUT(n1700), .C0(\adrram[1] ), .Z(n1711));
    PFUMX i1578 (.BLUT(n1670), .ALUT(n1671), .C0(\adrram[1] ), .Z(n1681));
    LUT4 i1656_3_lut (.A(\mem[12] [7]), .B(\mem[13] [7]), .C(\adrram[0] ), 
         .Z(n1759)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1656_3_lut.init = 16'hcaca;
    FD1P3AX mem_55__i0_i3 (.D(data[3]), .SP(we_N_63_enable_497), .CK(we_N_63), 
            .Q(\mem[55] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_55__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_55__i0_i2 (.D(data[2]), .SP(we_N_63_enable_497), .CK(we_N_63), 
            .Q(\mem[55] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_55__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_55__i0_i1 (.D(data[1]), .SP(we_N_63_enable_497), .CK(we_N_63), 
            .Q(\mem[55] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_55__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_54__i0_i7 (.D(data[7]), .SP(we_N_63_enable_505), .CK(we_N_63), 
            .Q(\mem[54] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_54__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_54__i0_i6 (.D(data[6]), .SP(we_N_63_enable_505), .CK(we_N_63), 
            .Q(\mem[54] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_54__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_43__i0_i3 (.D(data[3]), .SP(we_N_63_enable_511), .CK(we_N_63), 
            .Q(\mem[43] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_43__i0_i3.GSR = "ENABLED";
    PFUMX i1580 (.BLUT(n1674), .ALUT(n1675), .C0(\adrram[1] ), .Z(n1683));
    FD1P3AX mem_54__i0_i5 (.D(data[5]), .SP(we_N_63_enable_505), .CK(we_N_63), 
            .Q(\mem[54] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_54__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_54__i0_i4 (.D(data[4]), .SP(we_N_63_enable_505), .CK(we_N_63), 
            .Q(\mem[54] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_54__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_54__i0_i3 (.D(data[3]), .SP(we_N_63_enable_505), .CK(we_N_63), 
            .Q(\mem[54] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_54__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_54__i0_i2 (.D(data[2]), .SP(we_N_63_enable_505), .CK(we_N_63), 
            .Q(\mem[54] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_54__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_54__i0_i1 (.D(data[1]), .SP(we_N_63_enable_505), .CK(we_N_63), 
            .Q(\mem[54] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_54__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_43__i0_i2 (.D(data[2]), .SP(we_N_63_enable_511), .CK(we_N_63), 
            .Q(\mem[43] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_43__i0_i2.GSR = "ENABLED";
    PFUMX i1704 (.BLUT(n1798), .ALUT(n1799), .C0(\adrram[1] ), .Z(n1807));
    LUT4 i1787_3_lut (.A(\mem[58] [4]), .B(\mem[59] [4]), .C(\adrram[0] ), 
         .Z(n1890)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1787_3_lut.init = 16'hcaca;
    FD1P3AX mem_53__i0_i7 (.D(data[7]), .SP(we_N_63_enable_512), .CK(we_N_63), 
            .Q(\mem[53] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_53__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_53__i0_i6 (.D(data[6]), .SP(we_N_63_enable_512), .CK(we_N_63), 
            .Q(\mem[53] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_53__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_53__i0_i5 (.D(data[5]), .SP(we_N_63_enable_512), .CK(we_N_63), 
            .Q(\mem[53] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_53__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_53__i0_i4 (.D(data[4]), .SP(we_N_63_enable_512), .CK(we_N_63), 
            .Q(\mem[53] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_53__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_43__i0_i1 (.D(data[1]), .SP(we_N_63_enable_511), .CK(we_N_63), 
            .Q(\mem[43] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_43__i0_i1.GSR = "ENABLED";
    PFUMX i1828 (.BLUT(n1922), .ALUT(n1923), .C0(\adrram[1] ), .Z(n1931));
    PFUMX i1890 (.BLUT(n1984), .ALUT(n1985), .C0(\adrram[1] ), .Z(n1993));
    PFUMX i1455 (.BLUT(n1548), .ALUT(n1549), .C0(\adrram[1] ), .Z(n1558));
    LUT4 i1780_3_lut (.A(\mem[44] [4]), .B(\mem[45] [4]), .C(\adrram[0] ), 
         .Z(n1883)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1780_3_lut.init = 16'hcaca;
    LUT4 i1600_3_lut (.A(\mem[24] [5]), .B(\mem[25] [5]), .C(\adrram[0] ), 
         .Z(n1703)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1600_3_lut.init = 16'hcaca;
    LUT4 i1786_3_lut (.A(\mem[56] [4]), .B(\mem[57] [4]), .C(\adrram[0] ), 
         .Z(n1889)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1786_3_lut.init = 16'hcaca;
    LUT4 i1655_3_lut (.A(\mem[10] [7]), .B(\mem[11] [7]), .C(\adrram[0] ), 
         .Z(n1758)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1655_3_lut.init = 16'hcaca;
    LUT4 i1654_3_lut (.A(\mem[8] [7]), .B(\mem[9] [7]), .C(\adrram[0] ), 
         .Z(n1757)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1654_3_lut.init = 16'hcaca;
    LUT4 i1560_3_lut (.A(\mem[6] [4]), .B(\mem[7] [4]), .C(\adrram[0] ), 
         .Z(n1663)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1560_3_lut.init = 16'hcaca;
    LUT4 i1632_3_lut (.A(\mem[26] [6]), .B(\mem[27] [6]), .C(\adrram[0] ), 
         .Z(n1735)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1632_3_lut.init = 16'hcaca;
    LUT4 i1653_3_lut (.A(\mem[6] [7]), .B(\mem[7] [7]), .C(\adrram[0] ), 
         .Z(n1756)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1653_3_lut.init = 16'hcaca;
    LUT4 i1631_3_lut (.A(\mem[24] [6]), .B(\mem[25] [6]), .C(\adrram[0] ), 
         .Z(n1734)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1631_3_lut.init = 16'hcaca;
    LUT4 i1620_3_lut (.A(\mem[2] [6]), .B(\mem[3] [6]), .C(\adrram[0] ), 
         .Z(n1723)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1620_3_lut.init = 16'hcaca;
    LUT4 i1599_3_lut (.A(\mem[22] [5]), .B(\mem[23] [5]), .C(\adrram[0] ), 
         .Z(n1702)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1599_3_lut.init = 16'hcaca;
    LUT4 i1589_3_lut (.A(\mem[2] [5]), .B(\mem[3] [5]), .C(\adrram[0] ), 
         .Z(n1692)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1589_3_lut.init = 16'hcaca;
    LUT4 i1652_3_lut (.A(\mem[4] [7]), .B(\mem[5] [7]), .C(\adrram[0] ), 
         .Z(n1755)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1652_3_lut.init = 16'hcaca;
    LUT4 i1630_3_lut (.A(\mem[22] [6]), .B(\mem[23] [6]), .C(\adrram[0] ), 
         .Z(n1733)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1630_3_lut.init = 16'hcaca;
    LUT4 i1619_3_lut (.A(\mem[0] [6]), .B(\mem[1] [6]), .C(\adrram[0] ), 
         .Z(n1722)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1619_3_lut.init = 16'hcaca;
    PFUMX i1885 (.BLUT(n1974), .ALUT(n1975), .C0(\adrram[1] ), .Z(n1988));
    LUT4 i1598_3_lut (.A(\mem[20] [5]), .B(\mem[21] [5]), .C(\adrram[0] ), 
         .Z(n1701)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1598_3_lut.init = 16'hcaca;
    LUT4 i1588_3_lut (.A(\mem[0] [5]), .B(\mem[1] [5]), .C(\adrram[0] ), 
         .Z(n1691)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1588_3_lut.init = 16'hcaca;
    LUT4 i1559_3_lut (.A(\mem[4] [4]), .B(\mem[5] [4]), .C(\adrram[0] ), 
         .Z(n1662)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1559_3_lut.init = 16'hcaca;
    LUT4 i1629_3_lut (.A(\mem[20] [6]), .B(\mem[21] [6]), .C(\adrram[0] ), 
         .Z(n1732)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1629_3_lut.init = 16'hcaca;
    LUT4 i1651_3_lut (.A(\mem[2] [7]), .B(\mem[3] [7]), .C(\adrram[0] ), 
         .Z(n1754)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1651_3_lut.init = 16'hcaca;
    LUT4 i1650_3_lut (.A(\mem[0] [7]), .B(\mem[1] [7]), .C(\adrram[0] ), 
         .Z(n1753)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1650_3_lut.init = 16'hcaca;
    LUT4 i1475_3_lut (.A(\mem[22] [1]), .B(\mem[23] [1]), .C(\adrram[0] ), 
         .Z(n1578)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1475_3_lut.init = 16'hcaca;
    LUT4 i1785_3_lut (.A(\mem[54] [4]), .B(\mem[55] [4]), .C(\adrram[0] ), 
         .Z(n1888)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1785_3_lut.init = 16'hcaca;
    LUT4 i1903_3_lut (.A(\mem[42] [0]), .B(\mem[43] [0]), .C(\adrram[0] ), 
         .Z(n2006)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1903_3_lut.init = 16'hcaca;
    LUT4 i1784_3_lut (.A(\mem[52] [4]), .B(\mem[53] [4]), .C(\adrram[0] ), 
         .Z(n1887)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1784_3_lut.init = 16'hcaca;
    LUT4 i1779_3_lut (.A(\mem[42] [4]), .B(\mem[43] [4]), .C(\adrram[0] ), 
         .Z(n1882)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1779_3_lut.init = 16'hcaca;
    LUT4 i1597_3_lut (.A(\mem[18] [5]), .B(\mem[19] [5]), .C(\adrram[0] ), 
         .Z(n1700)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1597_3_lut.init = 16'hcaca;
    LUT4 i1566_3_lut (.A(\mem[18] [4]), .B(\mem[19] [4]), .C(\adrram[0] ), 
         .Z(n1669)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1566_3_lut.init = 16'hcaca;
    LUT4 i1558_3_lut (.A(\mem[2] [4]), .B(\mem[3] [4]), .C(\adrram[0] ), 
         .Z(n1661)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1558_3_lut.init = 16'hcaca;
    LUT4 i1474_3_lut (.A(\mem[20] [1]), .B(\mem[21] [1]), .C(\adrram[0] ), 
         .Z(n1577)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1474_3_lut.init = 16'hcaca;
    LUT4 i1902_3_lut (.A(\mem[40] [0]), .B(\mem[41] [0]), .C(\adrram[0] ), 
         .Z(n2005)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1902_3_lut.init = 16'hcaca;
    LUT4 i1628_3_lut (.A(\mem[18] [6]), .B(\mem[19] [6]), .C(\adrram[0] ), 
         .Z(n1731)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1628_3_lut.init = 16'hcaca;
    LUT4 i1778_3_lut (.A(\mem[40] [4]), .B(\mem[41] [4]), .C(\adrram[0] ), 
         .Z(n1881)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1778_3_lut.init = 16'hcaca;
    LUT4 i1596_3_lut (.A(\mem[16] [5]), .B(\mem[17] [5]), .C(\adrram[0] ), 
         .Z(n1699)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1596_3_lut.init = 16'hcaca;
    LUT4 i1565_3_lut (.A(\mem[16] [4]), .B(\mem[17] [4]), .C(\adrram[0] ), 
         .Z(n1668)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1565_3_lut.init = 16'hcaca;
    LUT4 i1557_3_lut (.A(\mem[0] [4]), .B(\mem[1] [4]), .C(\adrram[0] ), 
         .Z(n1660)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1557_3_lut.init = 16'hcaca;
    LUT4 i1469_3_lut (.A(\mem[10] [1]), .B(\mem[11] [1]), .C(\adrram[0] ), 
         .Z(n1572)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1469_3_lut.init = 16'hcaca;
    LUT4 i1527_3_lut (.A(\mem[2] [3]), .B(\mem[3] [3]), .C(\adrram[0] ), 
         .Z(n1630)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1527_3_lut.init = 16'hcaca;
    LUT4 i1526_3_lut (.A(\mem[0] [3]), .B(\mem[1] [3]), .C(\adrram[0] ), 
         .Z(n1629)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1526_3_lut.init = 16'hcaca;
    LUT4 i1880_3_lut (.A(\mem[58] [1]), .B(\mem[59] [1]), .C(\adrram[0] ), 
         .Z(n1983)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1880_3_lut.init = 16'hcaca;
    LUT4 i1815_3_lut (.A(\mem[52] [3]), .B(\mem[53] [3]), .C(\adrram[0] ), 
         .Z(n1918)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1815_3_lut.init = 16'hcaca;
    LUT4 i1816_3_lut (.A(\mem[54] [3]), .B(\mem[55] [3]), .C(\adrram[0] ), 
         .Z(n1919)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1816_3_lut.init = 16'hcaca;
    LUT4 i1687_3_lut (.A(\mem[44] [7]), .B(\mem[45] [7]), .C(\adrram[0] ), 
         .Z(n1790)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1687_3_lut.init = 16'hcaca;
    LUT4 i1688_3_lut (.A(\mem[46] [7]), .B(\mem[47] [7]), .C(\adrram[0] ), 
         .Z(n1791)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1688_3_lut.init = 16'hcaca;
    LUT4 i1689_3_lut (.A(\mem[48] [7]), .B(\mem[49] [7]), .C(\adrram[0] ), 
         .Z(n1792)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1689_3_lut.init = 16'hcaca;
    LUT4 i1690_3_lut (.A(\mem[50] [7]), .B(\mem[51] [7]), .C(\adrram[0] ), 
         .Z(n1793)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1690_3_lut.init = 16'hcaca;
    LUT4 i1817_3_lut (.A(\mem[56] [3]), .B(\mem[57] [3]), .C(\adrram[0] ), 
         .Z(n1920)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1817_3_lut.init = 16'hcaca;
    LUT4 i1818_3_lut (.A(\mem[58] [3]), .B(\mem[59] [3]), .C(\adrram[0] ), 
         .Z(n1921)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1818_3_lut.init = 16'hcaca;
    LUT4 i1691_3_lut (.A(\mem[52] [7]), .B(\mem[53] [7]), .C(\adrram[0] ), 
         .Z(n1794)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1691_3_lut.init = 16'hcaca;
    LUT4 i2272_2_lut_2_lut_3_lut_4_lut (.A(\adrram[1] ), .B(n2250), .C(n2248), 
         .D(\adrram[3] ), .Z(we_N_63_enable_231)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2272_2_lut_2_lut_3_lut_4_lut.init = 16'h0200;
    LUT4 i1692_3_lut (.A(\mem[54] [7]), .B(\mem[55] [7]), .C(\adrram[0] ), 
         .Z(n1795)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1692_3_lut.init = 16'hcaca;
    LUT4 i2182_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2257), .C(n2248), 
         .D(\adrram[3] ), .Z(we_N_63_enable_196)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2182_2_lut_2_lut_3_lut_4_lut.init = 16'h0002;
    LUT4 i1693_3_lut (.A(\mem[56] [7]), .B(\mem[57] [7]), .C(\adrram[0] ), 
         .Z(n1796)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1693_3_lut.init = 16'hcaca;
    LUT4 i1694_3_lut (.A(\mem[58] [7]), .B(\mem[59] [7]), .C(\adrram[0] ), 
         .Z(n1797)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1694_3_lut.init = 16'hcaca;
    LUT4 i1912_3_lut (.A(\mem[60] [0]), .B(\mem[61] [0]), .C(\adrram[0] ), 
         .Z(n2015)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1912_3_lut.init = 16'hcaca;
    LUT4 i1913_3_lut (.A(\mem[62] [0]), .B(\mem[63] [0]), .C(\adrram[0] ), 
         .Z(n2016)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1913_3_lut.init = 16'hcaca;
    LUT4 Select_638_i3_4_lut (.A(data_7__N_66[6]), .B(akku_o_c_6), .C(oe_N_57), 
         .D(n2247), .Z(data[6])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((D)+!B)) */ ;
    defparam Select_638_i3_4_lut.init = 16'ha0ec;
    LUT4 i1907_3_lut (.A(\mem[50] [0]), .B(\mem[51] [0]), .C(\adrram[0] ), 
         .Z(n2010)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1907_3_lut.init = 16'hcaca;
    LUT4 i2197_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2257), .C(n2249), 
         .D(\adrram[3] ), .Z(we_N_63_enable_343)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2197_2_lut_2_lut_3_lut_4_lut.init = 16'h0200;
    LUT4 i2216_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2257), .C(n2248), 
         .D(\adrram[3] ), .Z(we_N_63_enable_252)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2216_2_lut_2_lut_3_lut_4_lut.init = 16'h0200;
    LUT4 i2311_2_lut_2_lut_3_lut_4_lut (.A(\adrram[3] ), .B(n2249), .C(n2257), 
         .D(\adrram[2] ), .Z(we_N_63_enable_414)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2311_2_lut_2_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i2258_2_lut_2_lut_3_lut_4_lut (.A(\adrram[3] ), .B(n2249), .C(n2250), 
         .D(\adrram[1] ), .Z(we_N_63_enable_287)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2258_2_lut_2_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i2207_2_lut_2_lut_3_lut_4_lut (.A(\adrram[1] ), .B(n2259), .C(n2248), 
         .D(\adrram[3] ), .Z(we_N_63_enable_259)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i2207_2_lut_2_lut_3_lut_4_lut.init = 16'h0800;
    LUT4 i2288_2_lut_2_lut_3_lut_4_lut (.A(\adrram[1] ), .B(n2259), .C(n2249), 
         .D(\adrram[3] ), .Z(we_N_63_enable_376)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i2288_2_lut_2_lut_3_lut_4_lut.init = 16'h0008;
    LUT4 i2280_2_lut_2_lut_3_lut_4_lut (.A(\adrram[1] ), .B(n2259), .C(n2248), 
         .D(\adrram[3] ), .Z(we_N_63_enable_203)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i2280_2_lut_2_lut_3_lut_4_lut.init = 16'h0008;
    LUT4 i2269_2_lut_2_lut_3_lut_4_lut (.A(\adrram[1] ), .B(n2259), .C(n2249), 
         .D(\adrram[3] ), .Z(we_N_63_enable_350)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i2269_2_lut_2_lut_3_lut_4_lut.init = 16'h0800;
    LUT4 i1906_3_lut (.A(\mem[48] [0]), .B(\mem[49] [0]), .C(\adrram[0] ), 
         .Z(n2009)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1906_3_lut.init = 16'hcaca;
    LUT4 i2286_2_lut_2_lut_3_lut_4_lut (.A(\adrram[4] ), .B(n2258), .C(n2257), 
         .D(\adrram[2] ), .Z(we_N_63_enable_119)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2286_2_lut_2_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i2290_2_lut_2_lut_3_lut_4_lut (.A(\adrram[4] ), .B(n2258), .C(n2259), 
         .D(\adrram[1] ), .Z(we_N_63_enable_120)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2290_2_lut_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i2179_2_lut_2_lut_3_lut_4_lut (.A(\adrram[4] ), .B(n2258), .C(n2250), 
         .D(\adrram[1] ), .Z(we_N_63_enable_107)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2179_2_lut_2_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i2252_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2251), .C(n2249), 
         .D(\adrram[3] ), .Z(we_N_63_enable_301)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2252_2_lut_2_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i2314_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2251), .C(n2258), 
         .D(\adrram[4] ), .Z(we_N_63_enable_357)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2314_2_lut_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i2164_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2251), .C(n2248), 
         .D(\adrram[3] ), .Z(we_N_63_enable_210)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2164_2_lut_2_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i2360_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2251), .C(n2248), 
         .D(\adrram[3] ), .Z(we_N_63_enable_154)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2360_2_lut_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i2267_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2251), .C(n2249), 
         .D(\adrram[3] ), .Z(we_N_63_enable_266)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2267_2_lut_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i2249_2_lut_2_lut_3_lut_4_lut (.A(\adrram[1] ), .B(n2250), .C(n2249), 
         .D(\adrram[3] ), .Z(we_N_63_enable_308)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2249_2_lut_2_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i2357_2_lut_2_lut_3_lut_4_lut (.A(\adrram[1] ), .B(n2250), .C(n2248), 
         .D(\adrram[3] ), .Z(we_N_63_enable_161)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2357_2_lut_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i2167_2_lut_2_lut_3_lut_4_lut (.A(\adrram[1] ), .B(n2250), .C(n2258), 
         .D(\adrram[4] ), .Z(we_N_63_enable_144)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2167_2_lut_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i2264_2_lut_2_lut_3_lut_4_lut (.A(\adrram[1] ), .B(n2250), .C(n2249), 
         .D(\adrram[3] ), .Z(we_N_63_enable_273)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2264_2_lut_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i2278_2_lut_2_lut_3_lut_4_lut (.A(\adrram[1] ), .B(n2250), .C(n2248), 
         .D(\adrram[3] ), .Z(we_N_63_enable_217)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2278_2_lut_2_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i2188_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2251), .C(n2248), 
         .D(\adrram[3] ), .Z(we_N_63_enable_182)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2188_2_lut_2_lut_3_lut_4_lut.init = 16'h0002;
    LUT4 i2205_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2251), .C(n2258), 
         .D(\adrram[4] ), .Z(we_N_63_enable_117)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2205_2_lut_2_lut_3_lut_4_lut.init = 16'h0002;
    LUT4 i2255_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2251), .C(n2249), 
         .D(\adrram[3] ), .Z(we_N_63_enable_294)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2255_2_lut_2_lut_3_lut_4_lut.init = 16'h0002;
    LUT4 i2213_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2251), .C(n2249), 
         .D(\adrram[3] ), .Z(we_N_63_enable_329)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2213_2_lut_2_lut_3_lut_4_lut.init = 16'h0200;
    LUT4 i2225_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2251), .C(n2248), 
         .D(\adrram[3] ), .Z(we_N_63_enable_238)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2225_2_lut_2_lut_3_lut_4_lut.init = 16'h0200;
    LUT4 i2342_2_lut_2_lut_3_lut_4_lut (.A(\adrram[4] ), .B(n2255), .C(n2251), 
         .D(\adrram[2] ), .Z(we_N_63_enable_488)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i2342_2_lut_2_lut_3_lut_4_lut.init = 16'h0008;
    LUT4 i1136_2_lut_3_lut_4_lut (.A(\adrram[4] ), .B(n2255), .C(n2259), 
         .D(\adrram[1] ), .Z(we_N_63_enable_364)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1136_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i2348_2_lut_2_lut_3_lut_4_lut (.A(\adrram[4] ), .B(n2255), .C(n2250), 
         .D(\adrram[1] ), .Z(we_N_63_enable_461)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i2348_2_lut_2_lut_3_lut_4_lut.init = 16'h0800;
    LUT4 i2344_2_lut_2_lut_3_lut_4_lut (.A(\adrram[4] ), .B(n2255), .C(n2250), 
         .D(\adrram[1] ), .Z(we_N_63_enable_479)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i2344_2_lut_2_lut_3_lut_4_lut.init = 16'h0008;
    LUT4 i2350_2_lut_2_lut_3_lut_4_lut (.A(\adrram[4] ), .B(n2255), .C(n2251), 
         .D(\adrram[2] ), .Z(we_N_63_enable_452)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i2350_2_lut_2_lut_3_lut_4_lut.init = 16'h0800;
    LUT4 i2354_2_lut_2_lut_3_lut_4_lut (.A(\adrram[4] ), .B(n2255), .C(n2257), 
         .D(\adrram[2] ), .Z(we_N_63_enable_433)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i2354_2_lut_2_lut_3_lut_4_lut.init = 16'h0800;
    LUT4 i2173_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2257), .C(n2258), 
         .D(\adrram[4] ), .Z(we_N_63_enable_106)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2173_2_lut_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i2346_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2257), .C(n2255), 
         .D(\adrram[4] ), .Z(we_N_63_enable_470)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2346_2_lut_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i2194_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2257), .C(n2248), 
         .D(\adrram[3] ), .Z(we_N_63_enable_168)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2194_2_lut_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i2261_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2257), .C(n2249), 
         .D(\adrram[3] ), .Z(we_N_63_enable_280)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2261_2_lut_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i2246_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2257), .C(n2249), 
         .D(\adrram[3] ), .Z(we_N_63_enable_315)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2246_2_lut_2_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i2275_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2257), .C(n2248), 
         .D(\adrram[3] ), .Z(we_N_63_enable_224)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2275_2_lut_2_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i2293_2_lut_2_lut_3_lut_4_lut (.A(\adrram[4] ), .B(n2255), .C(n2251), 
         .D(\adrram[2] ), .Z(we_N_63_enable_121)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2293_2_lut_2_lut_3_lut_4_lut.init = 16'h0004;
    LUT4 i2296_2_lut_2_lut_3_lut_4_lut (.A(\adrram[4] ), .B(n2255), .C(n2250), 
         .D(\adrram[1] ), .Z(we_N_63_enable_122)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2296_2_lut_2_lut_3_lut_4_lut.init = 16'h0004;
    LUT4 i2320_2_lut_2_lut_3_lut_4_lut (.A(\adrram[4] ), .B(n2255), .C(n2251), 
         .D(\adrram[2] ), .Z(we_N_63_enable_475)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2320_2_lut_2_lut_3_lut_4_lut.init = 16'h0400;
    LUT4 i2202_2_lut_2_lut_3_lut_4_lut (.A(\adrram[4] ), .B(n2255), .C(n2259), 
         .D(\adrram[1] ), .Z(we_N_63_enable_416)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2202_2_lut_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 i2305_2_lut_2_lut_3_lut_4_lut (.A(\adrram[4] ), .B(n2255), .C(n2257), 
         .D(\adrram[2] ), .Z(we_N_63_enable_123)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2305_2_lut_2_lut_3_lut_4_lut.init = 16'h0004;
    LUT4 i2326_2_lut_2_lut_3_lut_4_lut (.A(\adrram[4] ), .B(n2255), .C(n2257), 
         .D(\adrram[2] ), .Z(we_N_63_enable_423)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2326_2_lut_2_lut_3_lut_4_lut.init = 16'h0400;
    LUT4 i2317_2_lut_2_lut_3_lut_4_lut (.A(\adrram[4] ), .B(n2255), .C(n2250), 
         .D(\adrram[1] ), .Z(we_N_63_enable_511)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2317_2_lut_2_lut_3_lut_4_lut.init = 16'h0400;
    LUT4 i2338_2_lut_2_lut_3_lut_4_lut (.A(\adrram[4] ), .B(n2258), .C(n2257), 
         .D(\adrram[2] ), .Z(we_N_63_enable_505)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2338_2_lut_2_lut_3_lut_4_lut.init = 16'h0200;
    LUT4 i2335_2_lut_2_lut_3_lut_4_lut (.A(\adrram[4] ), .B(n2258), .C(n2257), 
         .D(\adrram[2] ), .Z(we_N_63_enable_382)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2335_2_lut_2_lut_3_lut_4_lut.init = 16'h0002;
    LUT4 i2329_2_lut_2_lut_3_lut_4_lut (.A(\adrram[4] ), .B(n2258), .C(n2251), 
         .D(\adrram[2] ), .Z(we_N_63_enable_396)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2329_2_lut_2_lut_3_lut_4_lut.init = 16'h0002;
    LUT4 i2340_2_lut_2_lut_3_lut_4_lut (.A(\adrram[4] ), .B(n2258), .C(n2259), 
         .D(\adrram[1] ), .Z(we_N_63_enable_497)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2340_2_lut_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i1872_3_lut (.A(\mem[42] [1]), .B(\mem[43] [1]), .C(\adrram[0] ), 
         .Z(n1975)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1872_3_lut.init = 16'hcaca;
    LUT4 i2299_2_lut_2_lut_3_lut_4_lut (.A(\adrram[4] ), .B(n2258), .C(n2251), 
         .D(\adrram[2] ), .Z(we_N_63_enable_133)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2299_2_lut_2_lut_3_lut_4_lut.init = 16'h0200;
    LUT4 i2332_2_lut_2_lut_3_lut_4_lut (.A(\adrram[4] ), .B(n2258), .C(n2250), 
         .D(\adrram[1] ), .Z(we_N_63_enable_389)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2332_2_lut_2_lut_3_lut_4_lut.init = 16'h0002;
    LUT4 i2170_2_lut_2_lut_3_lut_4_lut (.A(\adrram[4] ), .B(n2258), .C(n2250), 
         .D(\adrram[1] ), .Z(we_N_63_enable_373)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2170_2_lut_2_lut_3_lut_4_lut.init = 16'h0200;
    LUT4 i2210_2_lut_2_lut_3_lut_4_lut (.A(\adrram[1] ), .B(n2259), .C(n2249), 
         .D(\adrram[3] ), .Z(we_N_63_enable_336)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2210_2_lut_2_lut_3_lut_4_lut.init = 16'h0400;
    LUT4 i637_1_lut (.A(\adrram[0] ), .Z(\pc_5__N_30[0] )) /* synthesis lut_function=(!(A)) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i637_1_lut.init = 16'h5555;
    LUT4 i1871_3_lut (.A(\mem[40] [1]), .B(\mem[41] [1]), .C(\adrram[0] ), 
         .Z(n1974)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1871_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_21 (.A(\adrram[0] ), .B(\adrram[1] ), .Z(n2251)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i1_2_lut_rep_21.init = 16'heeee;
    PFUMX i1918 (.BLUT(n2009), .ALUT(n2010), .C0(\adrram[1] ), .Z(n2021));
    LUT4 i1127_2_lut_rep_25 (.A(\adrram[5] ), .B(\adrram[3] ), .Z(n2255)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1127_2_lut_rep_25.init = 16'h8888;
    LUT4 i1_2_lut_rep_27 (.A(\adrram[0] ), .B(\adrram[1] ), .Z(n2257)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i1_2_lut_rep_27.init = 16'hbbbb;
    LUT4 i1_2_lut_rep_28 (.A(\adrram[3] ), .B(\adrram[5] ), .Z(n2258)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i1_2_lut_rep_28.init = 16'hbbbb;
    LUT4 i1446_3_lut (.A(\mem[26] [0]), .B(\mem[27] [0]), .C(\adrram[0] ), 
         .Z(n1549)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1446_3_lut.init = 16'hcaca;
    LUT4 i1129_2_lut_rep_29 (.A(\adrram[0] ), .B(\adrram[2] ), .Z(n2259)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1129_2_lut_rep_29.init = 16'h8888;
    LUT4 i1445_3_lut (.A(\mem[24] [0]), .B(\mem[25] [0]), .C(\adrram[0] ), 
         .Z(n1548)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1445_3_lut.init = 16'hcaca;
    LUT4 i1870_3_lut (.A(\mem[38] [1]), .B(\mem[39] [1]), .C(\adrram[0] ), 
         .Z(n1973)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1870_3_lut.init = 16'hcaca;
    LUT4 Select_643_i3_4_lut (.A(data_7__N_66[1]), .B(akku_o_c_1), .C(oe_N_57), 
         .D(n2247), .Z(data[1])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((D)+!B)) */ ;
    defparam Select_643_i3_4_lut.init = 16'ha0ec;
    LUT4 i1881_3_lut (.A(\mem[60] [1]), .B(\mem[61] [1]), .C(\adrram[0] ), 
         .Z(n1984)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1881_3_lut.init = 16'hcaca;
    LUT4 i1882_3_lut (.A(\mem[62] [1]), .B(\mem[63] [1]), .C(\adrram[0] ), 
         .Z(n1985)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1882_3_lut.init = 16'hcaca;
    LUT4 i1819_3_lut (.A(\mem[60] [3]), .B(\mem[61] [3]), .C(\adrram[0] ), 
         .Z(n1922)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1819_3_lut.init = 16'hcaca;
    LUT4 i1820_3_lut (.A(\mem[62] [3]), .B(\mem[63] [3]), .C(\adrram[0] ), 
         .Z(n1923)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1820_3_lut.init = 16'hcaca;
    LUT4 i1695_3_lut (.A(\mem[60] [7]), .B(\mem[61] [7]), .C(\adrram[0] ), 
         .Z(n1798)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1695_3_lut.init = 16'hcaca;
    LUT4 Select_639_i3_4_lut (.A(data_7__N_66[5]), .B(akku_o_c_5), .C(oe_N_57), 
         .D(n2247), .Z(data[5])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((D)+!B)) */ ;
    defparam Select_639_i3_4_lut.init = 16'ha0ec;
    LUT4 i1696_3_lut (.A(\mem[62] [7]), .B(\mem[63] [7]), .C(\adrram[0] ), 
         .Z(n1799)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1696_3_lut.init = 16'hcaca;
    LUT4 i1571_3_lut (.A(\mem[28] [4]), .B(\mem[29] [4]), .C(\adrram[0] ), 
         .Z(n1674)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1571_3_lut.init = 16'hcaca;
    LUT4 i1572_3_lut (.A(\mem[30] [4]), .B(\mem[31] [4]), .C(\adrram[0] ), 
         .Z(n1675)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1572_3_lut.init = 16'hcaca;
    LUT4 i1567_3_lut (.A(\mem[20] [4]), .B(\mem[21] [4]), .C(\adrram[0] ), 
         .Z(n1670)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1567_3_lut.init = 16'hcaca;
    LUT4 i1756_3_lut (.A(\mem[58] [5]), .B(\mem[59] [5]), .C(\adrram[0] ), 
         .Z(n1859)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1756_3_lut.init = 16'hcaca;
    LUT4 Select_640_i3_4_lut (.A(data_7__N_66[4]), .B(akku_o_c_4), .C(oe_N_57), 
         .D(n2247), .Z(data[4])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((D)+!B)) */ ;
    defparam Select_640_i3_4_lut.init = 16'ha0ec;
    LUT4 i1468_3_lut (.A(\mem[8] [1]), .B(\mem[9] [1]), .C(\adrram[0] ), 
         .Z(n1571)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1468_3_lut.init = 16'hcaca;
    LUT4 i1755_3_lut (.A(\mem[56] [5]), .B(\mem[57] [5]), .C(\adrram[0] ), 
         .Z(n1858)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1755_3_lut.init = 16'hcaca;
    LUT4 i1473_3_lut (.A(\mem[18] [1]), .B(\mem[19] [1]), .C(\adrram[0] ), 
         .Z(n1576)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1473_3_lut.init = 16'hcaca;
    LUT4 i1472_3_lut (.A(\mem[16] [1]), .B(\mem[17] [1]), .C(\adrram[0] ), 
         .Z(n1575)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1472_3_lut.init = 16'hcaca;
    LUT4 i1725_3_lut (.A(\mem[58] [6]), .B(\mem[59] [6]), .C(\adrram[0] ), 
         .Z(n1828)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1725_3_lut.init = 16'hcaca;
    LUT4 i1724_3_lut (.A(\mem[56] [6]), .B(\mem[57] [6]), .C(\adrram[0] ), 
         .Z(n1827)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1724_3_lut.init = 16'hcaca;
    LUT4 i1723_3_lut (.A(\mem[54] [6]), .B(\mem[55] [6]), .C(\adrram[0] ), 
         .Z(n1826)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1723_3_lut.init = 16'hcaca;
    LUT4 i1722_3_lut (.A(\mem[52] [6]), .B(\mem[53] [6]), .C(\adrram[0] ), 
         .Z(n1825)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1722_3_lut.init = 16'hcaca;
    LUT4 i1721_3_lut (.A(\mem[50] [6]), .B(\mem[51] [6]), .C(\adrram[0] ), 
         .Z(n1824)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1721_3_lut.init = 16'hcaca;
    LUT4 i1720_3_lut (.A(\mem[48] [6]), .B(\mem[49] [6]), .C(\adrram[0] ), 
         .Z(n1823)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1720_3_lut.init = 16'hcaca;
    LUT4 i2352_2_lut_2_lut_3_lut_4_lut (.A(\adrram[1] ), .B(n2259), .C(n2255), 
         .D(\adrram[4] ), .Z(we_N_63_enable_443)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2352_2_lut_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 Select_641_i3_4_lut (.A(data_7__N_66[3]), .B(akku_o_c_3), .C(oe_N_57), 
         .D(n2247), .Z(data[3])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((D)+!B)) */ ;
    defparam Select_641_i3_4_lut.init = 16'ha0ec;
    LUT4 i1570_3_lut (.A(\mem[26] [4]), .B(\mem[27] [4]), .C(\adrram[0] ), 
         .Z(n1673)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1570_3_lut.init = 16'hcaca;
    LUT4 i2308_2_lut_2_lut_3_lut_4_lut (.A(\adrram[1] ), .B(n2259), .C(n2249), 
         .D(\adrram[3] ), .Z(we_N_63_enable_407)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2308_2_lut_2_lut_3_lut_4_lut.init = 16'h0004;
    LUT4 i2323_2_lut_2_lut_3_lut_4_lut (.A(\adrram[1] ), .B(n2259), .C(n2255), 
         .D(\adrram[4] ), .Z(we_N_63_enable_446)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2323_2_lut_2_lut_3_lut_4_lut.init = 16'h0040;
    LUT4 i1569_3_lut (.A(\mem[24] [4]), .B(\mem[25] [4]), .C(\adrram[0] ), 
         .Z(n1672)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1569_3_lut.init = 16'hcaca;
    LUT4 i1869_3_lut (.A(\mem[36] [1]), .B(\mem[37] [1]), .C(\adrram[0] ), 
         .Z(n1972)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1869_3_lut.init = 16'hcaca;
    LUT4 i1719_3_lut (.A(\mem[46] [6]), .B(\mem[47] [6]), .C(\adrram[0] ), 
         .Z(n1822)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1719_3_lut.init = 16'hcaca;
    LUT4 i1718_3_lut (.A(\mem[44] [6]), .B(\mem[45] [6]), .C(\adrram[0] ), 
         .Z(n1821)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1718_3_lut.init = 16'hcaca;
    LUT4 i1717_3_lut (.A(\mem[42] [6]), .B(\mem[43] [6]), .C(\adrram[0] ), 
         .Z(n1820)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1717_3_lut.init = 16'hcaca;
    LUT4 i1754_3_lut (.A(\mem[54] [5]), .B(\mem[55] [5]), .C(\adrram[0] ), 
         .Z(n1857)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1754_3_lut.init = 16'hcaca;
    LUT4 i1753_3_lut (.A(\mem[52] [5]), .B(\mem[53] [5]), .C(\adrram[0] ), 
         .Z(n1856)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1753_3_lut.init = 16'hcaca;
    LUT4 i2185_2_lut_2_lut_3_lut_4_lut (.A(\adrram[1] ), .B(n2259), .C(n2248), 
         .D(\adrram[3] ), .Z(we_N_63_enable_189)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2185_2_lut_2_lut_3_lut_4_lut.init = 16'h0004;
    LUT4 i2283_2_lut_2_lut_3_lut_4_lut (.A(\adrram[1] ), .B(n2259), .C(n2258), 
         .D(\adrram[4] ), .Z(we_N_63_enable_118)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2283_2_lut_2_lut_3_lut_4_lut.init = 16'h0004;
    LUT4 i2219_2_lut_2_lut_3_lut_4_lut (.A(\adrram[1] ), .B(n2259), .C(n2248), 
         .D(\adrram[3] ), .Z(we_N_63_enable_245)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2219_2_lut_2_lut_3_lut_4_lut.init = 16'h0400;
    LUT4 i1849_3_lut (.A(\mem[58] [2]), .B(\mem[59] [2]), .C(\adrram[0] ), 
         .Z(n1952)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1849_3_lut.init = 16'hcaca;
    LUT4 i1848_3_lut (.A(\mem[56] [2]), .B(\mem[57] [2]), .C(\adrram[0] ), 
         .Z(n1951)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1848_3_lut.init = 16'hcaca;
    LUT4 i1467_3_lut (.A(\mem[6] [1]), .B(\mem[7] [1]), .C(\adrram[0] ), 
         .Z(n1570)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1467_3_lut.init = 16'hcaca;
    LUT4 i1471_3_lut (.A(\mem[14] [1]), .B(\mem[15] [1]), .C(\adrram[0] ), 
         .Z(n1574)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1471_3_lut.init = 16'hcaca;
    LUT4 i1466_3_lut (.A(\mem[4] [1]), .B(\mem[5] [1]), .C(\adrram[0] ), 
         .Z(n1569)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1466_3_lut.init = 16'hcaca;
    LUT4 i1750_3_lut (.A(\mem[46] [5]), .B(\mem[47] [5]), .C(\adrram[0] ), 
         .Z(n1853)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1750_3_lut.init = 16'hcaca;
    LUT4 i1749_3_lut (.A(\mem[44] [5]), .B(\mem[45] [5]), .C(\adrram[0] ), 
         .Z(n1852)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1749_3_lut.init = 16'hcaca;
    LUT4 i1564_3_lut (.A(\mem[14] [4]), .B(\mem[15] [4]), .C(\adrram[0] ), 
         .Z(n1667)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1564_3_lut.init = 16'hcaca;
    LUT4 i2302_2_lut_2_lut_3_lut_4_lut (.A(\adrram[1] ), .B(n2259), .C(n2258), 
         .D(\adrram[4] ), .Z(we_N_63_enable_512)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i2302_2_lut_2_lut_3_lut_4_lut.init = 16'h0400;
    LUT4 i1_2_lut_rep_18 (.A(\adrram[4] ), .B(\adrram[5] ), .Z(n2248)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i1_2_lut_rep_18.init = 16'heeee;
    LUT4 i1470_3_lut (.A(\mem[12] [1]), .B(\mem[13] [1]), .C(\adrram[0] ), 
         .Z(n1573)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1470_3_lut.init = 16'hcaca;
    LUT4 i1847_3_lut (.A(\mem[54] [2]), .B(\mem[55] [2]), .C(\adrram[0] ), 
         .Z(n1950)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1847_3_lut.init = 16'hcaca;
    LUT4 i1846_3_lut (.A(\mem[52] [2]), .B(\mem[53] [2]), .C(\adrram[0] ), 
         .Z(n1949)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1846_3_lut.init = 16'hcaca;
    LUT4 i1758_3_lut (.A(\mem[62] [5]), .B(\mem[63] [5]), .C(\adrram[0] ), 
         .Z(n1861)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1758_3_lut.init = 16'hcaca;
    LUT4 i1716_3_lut (.A(\mem[40] [6]), .B(\mem[41] [6]), .C(\adrram[0] ), 
         .Z(n1819)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1716_3_lut.init = 16'hcaca;
    LUT4 i1715_3_lut (.A(\mem[38] [6]), .B(\mem[39] [6]), .C(\adrram[0] ), 
         .Z(n1818)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1715_3_lut.init = 16'hcaca;
    LUT4 i1714_3_lut (.A(\mem[36] [6]), .B(\mem[37] [6]), .C(\adrram[0] ), 
         .Z(n1817)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1714_3_lut.init = 16'hcaca;
    LUT4 i1713_3_lut (.A(\mem[34] [6]), .B(\mem[35] [6]), .C(\adrram[0] ), 
         .Z(n1816)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1713_3_lut.init = 16'hcaca;
    LUT4 i1712_3_lut (.A(\mem[32] [6]), .B(\mem[33] [6]), .C(\adrram[0] ), 
         .Z(n1815)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1712_3_lut.init = 16'hcaca;
    LUT4 i1479_3_lut (.A(\mem[30] [1]), .B(\mem[31] [1]), .C(\adrram[0] ), 
         .Z(n1582)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1479_3_lut.init = 16'hcaca;
    LUT4 i1478_3_lut (.A(\mem[28] [1]), .B(\mem[29] [1]), .C(\adrram[0] ), 
         .Z(n1581)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1478_3_lut.init = 16'hcaca;
    LUT4 i1477_3_lut (.A(\mem[26] [1]), .B(\mem[27] [1]), .C(\adrram[0] ), 
         .Z(n1580)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1477_3_lut.init = 16'hcaca;
    LUT4 i1476_3_lut (.A(\mem[24] [1]), .B(\mem[25] [1]), .C(\adrram[0] ), 
         .Z(n1579)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1476_3_lut.init = 16'hcaca;
    LUT4 i1568_3_lut (.A(\mem[22] [4]), .B(\mem[23] [4]), .C(\adrram[0] ), 
         .Z(n1671)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1568_3_lut.init = 16'hcaca;
    LUT4 i1879_3_lut (.A(\mem[56] [1]), .B(\mem[57] [1]), .C(\adrram[0] ), 
         .Z(n1982)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1879_3_lut.init = 16'hcaca;
    LUT4 i1686_3_lut (.A(\mem[42] [7]), .B(\mem[43] [7]), .C(\adrram[0] ), 
         .Z(n1789)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1686_3_lut.init = 16'hcaca;
    LUT4 i1685_3_lut (.A(\mem[40] [7]), .B(\mem[41] [7]), .C(\adrram[0] ), 
         .Z(n1788)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1685_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_20 (.A(\adrram[2] ), .B(\adrram[0] ), .Z(n2250)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i1_2_lut_rep_20.init = 16'hbbbb;
    LUT4 i1684_3_lut (.A(\mem[38] [7]), .B(\mem[39] [7]), .C(\adrram[0] ), 
         .Z(n1787)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1684_3_lut.init = 16'hcaca;
    LUT4 i1683_3_lut (.A(\mem[36] [7]), .B(\mem[37] [7]), .C(\adrram[0] ), 
         .Z(n1786)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1683_3_lut.init = 16'hcaca;
    LUT4 i1814_3_lut (.A(\mem[50] [3]), .B(\mem[51] [3]), .C(\adrram[0] ), 
         .Z(n1917)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1814_3_lut.init = 16'hcaca;
    LUT4 i1813_3_lut (.A(\mem[48] [3]), .B(\mem[49] [3]), .C(\adrram[0] ), 
         .Z(n1916)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1813_3_lut.init = 16'hcaca;
    LUT4 i1682_3_lut (.A(\mem[34] [7]), .B(\mem[35] [7]), .C(\adrram[0] ), 
         .Z(n1785)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1682_3_lut.init = 16'hcaca;
    LUT4 i1681_3_lut (.A(\mem[32] [7]), .B(\mem[33] [7]), .C(\adrram[0] ), 
         .Z(n1784)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1681_3_lut.init = 16'hcaca;
    LUT4 i1812_3_lut (.A(\mem[46] [3]), .B(\mem[47] [3]), .C(\adrram[0] ), 
         .Z(n1915)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1812_3_lut.init = 16'hcaca;
    LUT4 i1811_3_lut (.A(\mem[44] [3]), .B(\mem[45] [3]), .C(\adrram[0] ), 
         .Z(n1914)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1811_3_lut.init = 16'hcaca;
    LUT4 i1878_3_lut (.A(\mem[54] [1]), .B(\mem[55] [1]), .C(\adrram[0] ), 
         .Z(n1981)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1878_3_lut.init = 16'hcaca;
    LUT4 i1877_3_lut (.A(\mem[52] [1]), .B(\mem[53] [1]), .C(\adrram[0] ), 
         .Z(n1980)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1877_3_lut.init = 16'hcaca;
    LUT4 i1911_3_lut (.A(\mem[58] [0]), .B(\mem[59] [0]), .C(\adrram[0] ), 
         .Z(n2014)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1911_3_lut.init = 16'hcaca;
    LUT4 i1910_3_lut (.A(\mem[56] [0]), .B(\mem[57] [0]), .C(\adrram[0] ), 
         .Z(n2013)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1910_3_lut.init = 16'hcaca;
    LUT4 i1810_3_lut (.A(\mem[42] [3]), .B(\mem[43] [3]), .C(\adrram[0] ), 
         .Z(n1913)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1810_3_lut.init = 16'hcaca;
    LUT4 i1809_3_lut (.A(\mem[40] [3]), .B(\mem[41] [3]), .C(\adrram[0] ), 
         .Z(n1912)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1809_3_lut.init = 16'hcaca;
    LUT4 i1808_3_lut (.A(\mem[38] [3]), .B(\mem[39] [3]), .C(\adrram[0] ), 
         .Z(n1911)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1808_3_lut.init = 16'hcaca;
    LUT4 i1807_3_lut (.A(\mem[36] [3]), .B(\mem[37] [3]), .C(\adrram[0] ), 
         .Z(n1910)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1807_3_lut.init = 16'hcaca;
    LUT4 i1876_3_lut (.A(\mem[50] [1]), .B(\mem[51] [1]), .C(\adrram[0] ), 
         .Z(n1979)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1876_3_lut.init = 16'hcaca;
    PFUMX i1921 (.BLUT(n2015), .ALUT(n2016), .C0(\adrram[1] ), .Z(n2024));
    LUT4 i1875_3_lut (.A(\mem[48] [1]), .B(\mem[49] [1]), .C(\adrram[0] ), 
         .Z(n1978)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1875_3_lut.init = 16'hcaca;
    LUT4 i1806_3_lut (.A(\mem[34] [3]), .B(\mem[35] [3]), .C(\adrram[0] ), 
         .Z(n1909)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1806_3_lut.init = 16'hcaca;
    LUT4 i1805_3_lut (.A(\mem[32] [3]), .B(\mem[33] [3]), .C(\adrram[0] ), 
         .Z(n1908)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1805_3_lut.init = 16'hcaca;
    LUT4 i1510_3_lut (.A(\mem[30] [2]), .B(\mem[31] [2]), .C(\adrram[0] ), 
         .Z(n1613)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1510_3_lut.init = 16'hcaca;
    LUT4 i1509_3_lut (.A(\mem[28] [2]), .B(\mem[29] [2]), .C(\adrram[0] ), 
         .Z(n1612)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1509_3_lut.init = 16'hcaca;
    LUT4 i1508_3_lut (.A(\mem[26] [2]), .B(\mem[27] [2]), .C(\adrram[0] ), 
         .Z(n1611)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1508_3_lut.init = 16'hcaca;
    PFUMX i1703 (.BLUT(n1796), .ALUT(n1797), .C0(\adrram[1] ), .Z(n1806));
    LUT4 i1909_3_lut (.A(\mem[54] [0]), .B(\mem[55] [0]), .C(\adrram[0] ), 
         .Z(n2012)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1909_3_lut.init = 16'hcaca;
    LUT4 i1873_3_lut (.A(\mem[44] [1]), .B(\mem[45] [1]), .C(\adrram[0] ), 
         .Z(n1976)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1873_3_lut.init = 16'hcaca;
    LUT4 i1874_3_lut (.A(\mem[46] [1]), .B(\mem[47] [1]), .C(\adrram[0] ), 
         .Z(n1977)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1874_3_lut.init = 16'hcaca;
    LUT4 i1908_3_lut (.A(\mem[52] [0]), .B(\mem[53] [0]), .C(\adrram[0] ), 
         .Z(n2011)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1908_3_lut.init = 16'hcaca;
    LUT4 i1507_3_lut (.A(\mem[24] [2]), .B(\mem[25] [2]), .C(\adrram[0] ), 
         .Z(n1610)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1507_3_lut.init = 16'hcaca;
    LUT4 i1506_3_lut (.A(\mem[22] [2]), .B(\mem[23] [2]), .C(\adrram[0] ), 
         .Z(n1609)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1506_3_lut.init = 16'hcaca;
    FD1P3AX mem_53__i0_i3 (.D(data[3]), .SP(we_N_63_enable_512), .CK(we_N_63), 
            .Q(\mem[53] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(66[9] 75[16])
    defparam mem_53__i0_i3.GSR = "ENABLED";
    LUT4 i1444_3_lut (.A(\mem[22] [0]), .B(\mem[23] [0]), .C(\adrram[0] ), 
         .Z(n1547)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1444_3_lut.init = 16'hcaca;
    LUT4 i1443_3_lut (.A(\mem[20] [0]), .B(\mem[21] [0]), .C(\adrram[0] ), 
         .Z(n1546)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1443_3_lut.init = 16'hcaca;
    LUT4 i1502_3_lut (.A(\mem[14] [2]), .B(\mem[15] [2]), .C(\adrram[0] ), 
         .Z(n1605)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1502_3_lut.init = 16'hcaca;
    PFUMX i1702 (.BLUT(n1794), .ALUT(n1795), .C0(\adrram[1] ), .Z(n1805));
    LUT4 i1503_3_lut (.A(\mem[16] [2]), .B(\mem[17] [2]), .C(\adrram[0] ), 
         .Z(n1606)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1503_3_lut.init = 16'hcaca;
    PFUMX i1827 (.BLUT(n1920), .ALUT(n1921), .C0(\adrram[1] ), .Z(n1930));
    PFUMX i1701 (.BLUT(n1792), .ALUT(n1793), .C0(\adrram[1] ), .Z(n1804));
    PFUMX i1700 (.BLUT(n1790), .ALUT(n1791), .C0(\adrram[1] ), .Z(n1803));
    PFUMX i1826 (.BLUT(n1918), .ALUT(n1919), .C0(\adrram[1] ), .Z(n1929));
    PFUMX i1485 (.BLUT(n1577), .ALUT(n1578), .C0(\adrram[1] ), .Z(n1588));
    PFUMX i1916 (.BLUT(n2005), .ALUT(n2006), .C0(\adrram[1] ), .Z(n2019));
    PFUMX i1795 (.BLUT(n1887), .ALUT(n1888), .C0(\adrram[1] ), .Z(n1898));
    PFUMX i1666 (.BLUT(n1753), .ALUT(n1754), .C0(\adrram[1] ), .Z(n1769));
    PFUMX i1763 (.BLUT(n1854), .ALUT(n1855), .C0(\adrram[1] ), .Z(n1866));
    PFUMX i1574 (.BLUT(n1662), .ALUT(n1663), .C0(\adrram[1] ), .Z(n1677));
    PFUMX i1604 (.BLUT(n1691), .ALUT(n1692), .C0(\adrram[1] ), .Z(n1707));
    PFUMX i1609 (.BLUT(n1701), .ALUT(n1702), .C0(\adrram[1] ), .Z(n1712));
    PFUMX i1635 (.BLUT(n1722), .ALUT(n1723), .C0(\adrram[1] ), .Z(n1738));
    PFUMX i1640 (.BLUT(n1732), .ALUT(n1733), .C0(\adrram[1] ), .Z(n1743));
    PFUMX i1859 (.BLUT(n1953), .ALUT(n1954), .C0(\adrram[1] ), .Z(n1962));
    PFUMX i1667 (.BLUT(n1755), .ALUT(n1756), .C0(\adrram[1] ), .Z(n1770));
    PFUMX i1641 (.BLUT(n1734), .ALUT(n1735), .C0(\adrram[1] ), .Z(n1744));
    PFUMX i1668 (.BLUT(n1757), .ALUT(n1758), .C0(\adrram[1] ), .Z(n1771));
    PFUMX i1605 (.BLUT(n1693), .ALUT(n1694), .C0(\adrram[1] ), .Z(n1708));
    PFUMX i1610 (.BLUT(n1703), .ALUT(n1704), .C0(\adrram[1] ), .Z(n1713));
    PFUMX i1793 (.BLUT(n1883), .ALUT(n1884), .C0(\adrram[1] ), .Z(n1896));
    PFUMX i1796 (.BLUT(n1889), .ALUT(n1890), .C0(\adrram[1] ), .Z(n1899));
    PFUMX i1669 (.BLUT(n1759), .ALUT(n1760), .C0(\adrram[1] ), .Z(n1772));
    PFUMX i1642 (.BLUT(n1736), .ALUT(n1737), .C0(\adrram[1] ), .Z(n1745));
    PFUMX i1670 (.BLUT(n1761), .ALUT(n1762), .C0(\adrram[1] ), .Z(n1773));
    PFUMX i1636 (.BLUT(n1724), .ALUT(n1725), .C0(\adrram[1] ), .Z(n1739));
    PFUMX i1797 (.BLUT(n1891), .ALUT(n1892), .C0(\adrram[1] ), .Z(n1900));
    PFUMX i1611 (.BLUT(n1705), .ALUT(n1706), .C0(\adrram[1] ), .Z(n1714));
    PFUMX i1671 (.BLUT(n1763), .ALUT(n1764), .C0(\adrram[1] ), .Z(n1774));
    PFUMX i1914 (.BLUT(n2001), .ALUT(n2002), .C0(\adrram[1] ), .Z(n2017));
    PFUMX i1672 (.BLUT(n1765), .ALUT(n1766), .C0(\adrram[1] ), .Z(n1775));
    PFUMX i1543 (.BLUT(n1631), .ALUT(n1632), .C0(\adrram[1] ), .Z(n1646));
    PFUMX i1575 (.BLUT(n1664), .ALUT(n1665), .C0(\adrram[1] ), .Z(n1678));
    PFUMX i1637 (.BLUT(n1726), .ALUT(n1727), .C0(\adrram[1] ), .Z(n1740));
    PFUMX i1456 (.BLUT(n1550), .ALUT(n1551), .C0(\adrram[1] ), .Z(n1559));
    LUT4 i1501_3_lut (.A(\mem[12] [2]), .B(\mem[13] [2]), .C(\adrram[0] ), 
         .Z(n1604)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1501_3_lut.init = 16'hcaca;
    PFUMX i1606 (.BLUT(n1695), .ALUT(n1696), .C0(\adrram[1] ), .Z(n1709));
    PFUMX i1766 (.BLUT(n1860), .ALUT(n1861), .C0(\adrram[1] ), .Z(n1869));
    PFUMX i1790 (.BLUT(n1877), .ALUT(n1878), .C0(\adrram[1] ), .Z(n1893));
    PFUMX i1673 (.BLUT(n1767), .ALUT(n1768), .C0(\adrram[1] ), .Z(n1776));
    LUT4 i1500_3_lut (.A(\mem[10] [2]), .B(\mem[11] [2]), .C(\adrram[0] ), 
         .Z(n1603)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1500_3_lut.init = 16'hcaca;
    PFUMX i1576 (.BLUT(n1666), .ALUT(n1667), .C0(\adrram[1] ), .Z(n1679));
    PFUMX i1794 (.BLUT(n1885), .ALUT(n1886), .C0(\adrram[1] ), .Z(n1897));
    PFUMX i1449 (.BLUT(n1536), .ALUT(n1537), .C0(\adrram[1] ), .Z(n1552));
    LUT4 i1499_3_lut (.A(\mem[8] [2]), .B(\mem[9] [2]), .C(\adrram[0] ), 
         .Z(n1602)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1499_3_lut.init = 16'hcaca;
    PFUMX i1607 (.BLUT(n1697), .ALUT(n1698), .C0(\adrram[1] ), .Z(n1710));
    LUT4 i1498_3_lut (.A(\mem[6] [2]), .B(\mem[7] [2]), .C(\adrram[0] ), 
         .Z(n1601)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1498_3_lut.init = 16'hcaca;
    PFUMX i1791 (.BLUT(n1879), .ALUT(n1880), .C0(\adrram[1] ), .Z(n1894));
    PFUMX i1883 (.BLUT(n1970), .ALUT(n1971), .C0(\adrram[1] ), .Z(n1986));
    LUT4 i1497_3_lut (.A(\mem[4] [2]), .B(\mem[5] [2]), .C(\adrram[0] ), 
         .Z(n1600)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1497_3_lut.init = 16'hcaca;
    PFUMX i1638 (.BLUT(n1728), .ALUT(n1729), .C0(\adrram[1] ), .Z(n1741));
    PFUMX i1915 (.BLUT(n2003), .ALUT(n2004), .C0(\adrram[1] ), .Z(n2018));
    LUT4 i1496_3_lut (.A(\mem[2] [2]), .B(\mem[3] [2]), .C(\adrram[0] ), 
         .Z(n1599)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1496_3_lut.init = 16'hcaca;
    PFUMX i1917 (.BLUT(n2007), .ALUT(n2008), .C0(\adrram[1] ), .Z(n2020));
    LUT4 i1495_3_lut (.A(\mem[0] [2]), .B(\mem[1] [2]), .C(\adrram[0] ), 
         .Z(n1598)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1495_3_lut.init = 16'hcaca;
    PFUMX i1792 (.BLUT(n1881), .ALUT(n1882), .C0(\adrram[1] ), .Z(n1895));
    PFUMX i1639 (.BLUT(n1730), .ALUT(n1731), .C0(\adrram[1] ), .Z(n1742));
    PFUMX i1450 (.BLUT(n1538), .ALUT(n1539), .C0(\adrram[1] ), .Z(n1553));
    LUT4 i1_2_lut_rep_19 (.A(\adrram[5] ), .B(\adrram[4] ), .Z(n2249)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/70735/desktop/cpu_l/sram64kx8_lcm.vhd(73[21:47])
    defparam i1_2_lut_rep_19.init = 16'hbbbb;
    LUT4 i1928_3_lut (.A(n2029), .B(n2030), .C(\adrram[4] ), .Z(n2031)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1928_3_lut.init = 16'hcaca;
    PFUMX i1884 (.BLUT(n1972), .ALUT(n1973), .C0(\adrram[1] ), .Z(n1987));
    PFUMX i1735 (.BLUT(n1829), .ALUT(n1830), .C0(\adrram[1] ), .Z(n1838));
    PFUMX i1544 (.BLUT(n1633), .ALUT(n1634), .C0(\adrram[1] ), .Z(n1647));
    PFUMX i1545 (.BLUT(n1635), .ALUT(n1636), .C0(\adrram[1] ), .Z(n1648));
    PFUMX i1546 (.BLUT(n1637), .ALUT(n1638), .C0(\adrram[1] ), .Z(n1649));
    PFUMX i1547 (.BLUT(n1639), .ALUT(n1640), .C0(\adrram[1] ), .Z(n1650));
    PFUMX i1548 (.BLUT(n1641), .ALUT(n1642), .C0(\adrram[1] ), .Z(n1651));
    PFUMX i1549 (.BLUT(n1643), .ALUT(n1644), .C0(\adrram[1] ), .Z(n1652));
    PFUMX i1451 (.BLUT(n1540), .ALUT(n1541), .C0(\adrram[1] ), .Z(n1554));
    PFUMX i1452 (.BLUT(n1542), .ALUT(n1543), .C0(\adrram[1] ), .Z(n1555));
    PFUMX i1852 (.BLUT(n1939), .ALUT(n1940), .C0(\adrram[1] ), .Z(n1955));
    PFUMX i1853 (.BLUT(n1941), .ALUT(n1942), .C0(\adrram[1] ), .Z(n1956));
    PFUMX i1453 (.BLUT(n1544), .ALUT(n1545), .C0(\adrram[1] ), .Z(n1556));
    PFUMX i1854 (.BLUT(n1943), .ALUT(n1944), .C0(\adrram[1] ), .Z(n1957));
    PFUMX i1855 (.BLUT(n1945), .ALUT(n1946), .C0(\adrram[1] ), .Z(n1958));
    PFUMX i1759 (.BLUT(n1846), .ALUT(n1847), .C0(\adrram[1] ), .Z(n1862));
    PFUMX i1856 (.BLUT(n1947), .ALUT(n1948), .C0(\adrram[1] ), .Z(n1959));
    PFUMX i1760 (.BLUT(n1848), .ALUT(n1849), .C0(\adrram[1] ), .Z(n1863));
    PFUMX i1761 (.BLUT(n1850), .ALUT(n1851), .C0(\adrram[1] ), .Z(n1864));
    PFUMX i1480 (.BLUT(n1567), .ALUT(n1568), .C0(\adrram[1] ), .Z(n1583));
    LUT4 i1463_3_lut (.A(n1564), .B(n1565), .C(\adrram[4] ), .Z(n1566)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1463_3_lut.init = 16'hcaca;
    LUT4 i1897_3_lut (.A(n1998), .B(n1999), .C(\adrram[4] ), .Z(n2000)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1897_3_lut.init = 16'hcaca;
    LUT4 i1494_3_lut (.A(n1595), .B(n1596), .C(\adrram[4] ), .Z(n1597)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1494_3_lut.init = 16'hcaca;
    LUT4 i1866_3_lut (.A(n1967), .B(n1968), .C(\adrram[4] ), .Z(n1969)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1866_3_lut.init = 16'hcaca;
    LUT4 i1525_3_lut (.A(n1626), .B(n1627), .C(\adrram[4] ), .Z(n1628)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1525_3_lut.init = 16'hcaca;
    LUT4 i1835_3_lut (.A(n1936), .B(n1937), .C(\adrram[4] ), .Z(n1938)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1835_3_lut.init = 16'hcaca;
    LUT4 i1556_3_lut (.A(n1657), .B(n1658), .C(\adrram[4] ), .Z(n1659)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1556_3_lut.init = 16'hcaca;
    LUT4 i1804_3_lut (.A(n1905), .B(n1906), .C(\adrram[4] ), .Z(n1907)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1804_3_lut.init = 16'hcaca;
    LUT4 i1587_3_lut (.A(n1688), .B(n1689), .C(\adrram[4] ), .Z(n1690)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1587_3_lut.init = 16'hcaca;
    LUT4 i1773_3_lut (.A(n1874), .B(n1875), .C(\adrram[4] ), .Z(n1876)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1773_3_lut.init = 16'hcaca;
    LUT4 i1618_3_lut (.A(n1719), .B(n1720), .C(\adrram[4] ), .Z(n1721)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1618_3_lut.init = 16'hcaca;
    LUT4 i1742_3_lut (.A(n1843), .B(n1844), .C(\adrram[4] ), .Z(n1845)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1742_3_lut.init = 16'hcaca;
    LUT4 i1649_3_lut (.A(n1750), .B(n1751), .C(\adrram[4] ), .Z(n1752)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1649_3_lut.init = 16'hcaca;
    LUT4 i1711_3_lut (.A(n1812), .B(n1813), .C(\adrram[4] ), .Z(n1814)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1711_3_lut.init = 16'hcaca;
    LUT4 i1680_3_lut (.A(n1781), .B(n1782), .C(\adrram[4] ), .Z(n1783)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1680_3_lut.init = 16'hcaca;
    LUT4 i1505_3_lut (.A(\mem[20] [2]), .B(\mem[21] [2]), .C(\adrram[0] ), 
         .Z(n1608)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1505_3_lut.init = 16'hcaca;
    LUT4 i1504_3_lut (.A(\mem[18] [2]), .B(\mem[19] [2]), .C(\adrram[0] ), 
         .Z(n1607)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1504_3_lut.init = 16'hcaca;
    
endmodule
//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

