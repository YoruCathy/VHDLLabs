// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.10.0.111.2
// Netlist written on Wed Dec 09 16:38:54 2020
//
// Verilog Description of module cpu2system
//

module cpu2system (clk, reset, akku_o, disp2);   // c:/users/70735/desktop/cpu/cpu2system.vhd(8[8:18])
    input clk;   // c:/users/70735/desktop/cpu/cpu2system.vhd(9[13:16])
    input reset;   // c:/users/70735/desktop/cpu/cpu2system.vhd(10[13:18])
    output [8:0]akku_o;   // c:/users/70735/desktop/cpu/cpu2system.vhd(11[13:19])
    output [8:0]disp2;   // c:/users/70735/desktop/cpu/cpu2system.vhd(12[4:9])
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/70735/desktop/cpu/cpu2system.vhd(9[13:16])
    wire we_N_63 /* synthesis is_clock=1, is_inv_clock=1, SET_AS_NETWORK=\CPU/we_N_63 */ ;   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(13[13:15])
    
    wire GND_net, reset_c, akku_o_c_8, akku_o_c_7, akku_o_c_6, akku_o_c_5, 
        akku_o_c_4, akku_o_c_3, akku_o_c_2, akku_o_c_1, akku_o_c_0;
    wire [7:0]data;   // c:/users/70735/desktop/cpu/cpu2system.vhd(39[13:17])
    wire [15:0]adrram;   // c:/users/70735/desktop/cpu/cpu2system.vhd(40[13:19])
    wire [5:0]pc_5__N_30;
    
    wire oe_N_57, n2310, n2306, n2305, VCC_net, we_N_63_enable_315, 
        we_N_63_enable_259, n2314, n2313, we_N_63_enable_187;
    
    VHI i2444 (.Z(VCC_net));
    OB disp2_pad_2 (.I(GND_net), .O(disp2[2]));   // c:/users/70735/desktop/cpu/cpu2system.vhd(12[4:9])
    OB disp2_pad_3 (.I(GND_net), .O(disp2[3]));   // c:/users/70735/desktop/cpu/cpu2system.vhd(12[4:9])
    OB disp2_pad_4 (.I(GND_net), .O(disp2[4]));   // c:/users/70735/desktop/cpu/cpu2system.vhd(12[4:9])
    OB disp2_pad_5 (.I(GND_net), .O(disp2[5]));   // c:/users/70735/desktop/cpu/cpu2system.vhd(12[4:9])
    OB disp2_pad_6 (.I(GND_net), .O(disp2[6]));   // c:/users/70735/desktop/cpu/cpu2system.vhd(12[4:9])
    OB disp2_pad_7 (.I(GND_net), .O(disp2[7]));   // c:/users/70735/desktop/cpu/cpu2system.vhd(12[4:9])
    OB disp2_pad_8 (.I(GND_net), .O(disp2[8]));   // c:/users/70735/desktop/cpu/cpu2system.vhd(12[4:9])
    OB akku_o_pad_0 (.I(akku_o_c_0), .O(akku_o[0]));   // c:/users/70735/desktop/cpu/cpu2system.vhd(11[13:19])
    OB akku_o_pad_1 (.I(akku_o_c_1), .O(akku_o[1]));   // c:/users/70735/desktop/cpu/cpu2system.vhd(11[13:19])
    OB akku_o_pad_2 (.I(akku_o_c_2), .O(akku_o[2]));   // c:/users/70735/desktop/cpu/cpu2system.vhd(11[13:19])
    OB akku_o_pad_3 (.I(akku_o_c_3), .O(akku_o[3]));   // c:/users/70735/desktop/cpu/cpu2system.vhd(11[13:19])
    OB akku_o_pad_4 (.I(akku_o_c_4), .O(akku_o[4]));   // c:/users/70735/desktop/cpu/cpu2system.vhd(11[13:19])
    OB akku_o_pad_5 (.I(akku_o_c_5), .O(akku_o[5]));   // c:/users/70735/desktop/cpu/cpu2system.vhd(11[13:19])
    OB akku_o_pad_6 (.I(akku_o_c_6), .O(akku_o[6]));   // c:/users/70735/desktop/cpu/cpu2system.vhd(11[13:19])
    OB akku_o_pad_7 (.I(akku_o_c_7), .O(akku_o[7]));   // c:/users/70735/desktop/cpu/cpu2system.vhd(11[13:19])
    OB akku_o_pad_8 (.I(akku_o_c_8), .O(akku_o[8]));   // c:/users/70735/desktop/cpu/cpu2system.vhd(11[13:19])
    IB reset_pad (.I(reset), .O(reset_c));   // c:/users/70735/desktop/cpu/cpu2system.vhd(10[13:18])
    IB clk_pad (.I(clk), .O(clk_c));   // c:/users/70735/desktop/cpu/cpu2system.vhd(9[13:16])
    OB disp2_pad_0 (.I(GND_net), .O(disp2[0]));   // c:/users/70735/desktop/cpu/cpu2system.vhd(12[4:9])
    OB disp2_pad_1 (.I(GND_net), .O(disp2[1]));   // c:/users/70735/desktop/cpu/cpu2system.vhd(12[4:9])
    VLO i1 (.Z(GND_net));
    CPU8BIT2 CPU (.\adrram[0] (adrram[0]), .clk_c(clk_c), .akku_o_c_0(akku_o_c_0), 
            .pc_5__N_30({Open_0, Open_1, Open_2, Open_3, Open_4, pc_5__N_30[0]}), 
            .data({data}), .akku_o_c_8(akku_o_c_8), .akku_o_c_7(akku_o_c_7), 
            .akku_o_c_6(akku_o_c_6), .akku_o_c_5(akku_o_c_5), .akku_o_c_4(akku_o_c_4), 
            .akku_o_c_3(akku_o_c_3), .akku_o_c_2(akku_o_c_2), .akku_o_c_1(akku_o_c_1), 
            .\adrram[5] (adrram[5]), .\adrram[4] (adrram[4]), .\adrram[3] (adrram[3]), 
            .\adrram[2] (adrram[2]), .\adrram[1] (adrram[1]), .n2313(n2313), 
            .n2310(n2310), .we_N_63_enable_259(we_N_63_enable_259), .n2314(n2314), 
            .we_N_63_enable_315(we_N_63_enable_315), .n2306(n2306), .we_N_63_enable_187(we_N_63_enable_187), 
            .reset_c(reset_c), .we_N_63(we_N_63), .oe_N_57(oe_N_57), .n2305(n2305), 
            .GND_net(GND_net));   // c:/users/70735/desktop/cpu/cpu2system.vhd(46[10:18])
    TSALL TSALL_INST (.TSALL(GND_net));
    GSR GSR_INST (.GSR(reset_c));
    sram64kx8 RAM (.we_N_63(we_N_63), .data({data}), .we_N_63_enable_315(we_N_63_enable_315), 
            .we_N_63_enable_259(we_N_63_enable_259), .we_N_63_enable_187(we_N_63_enable_187), 
            .akku_o_c_0(akku_o_c_0), .oe_N_57(oe_N_57), .n2305(n2305), 
            .akku_o_c_5(akku_o_c_5), .\adrram[0] (adrram[0]), .\adrram[2] (adrram[2]), 
            .n2314(n2314), .\adrram[5] (adrram[5]), .\adrram[3] (adrram[3]), 
            .\adrram[1] (adrram[1]), .n2306(n2306), .n2310(n2310), .akku_o_c_4(akku_o_c_4), 
            .akku_o_c_3(akku_o_c_3), .n2313(n2313), .\pc_5__N_30[0] (pc_5__N_30[0]), 
            .\adrram[4] (adrram[4]), .akku_o_c_6(akku_o_c_6), .akku_o_c_2(akku_o_c_2), 
            .akku_o_c_1(akku_o_c_1), .akku_o_c_7(akku_o_c_7));   // c:/users/70735/desktop/cpu/cpu2system.vhd(47[10:19])
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    
endmodule
//
// Verilog Description of module CPU8BIT2
//

module CPU8BIT2 (\adrram[0] , clk_c, akku_o_c_0, pc_5__N_30, data, 
            akku_o_c_8, akku_o_c_7, akku_o_c_6, akku_o_c_5, akku_o_c_4, 
            akku_o_c_3, akku_o_c_2, akku_o_c_1, \adrram[5] , \adrram[4] , 
            \adrram[3] , \adrram[2] , \adrram[1] , n2313, n2310, we_N_63_enable_259, 
            n2314, we_N_63_enable_315, n2306, we_N_63_enable_187, reset_c, 
            we_N_63, oe_N_57, n2305, GND_net);
    output \adrram[0] ;
    input clk_c;
    output akku_o_c_0;
    input [5:0]pc_5__N_30;
    input [7:0]data;
    output akku_o_c_8;
    output akku_o_c_7;
    output akku_o_c_6;
    output akku_o_c_5;
    output akku_o_c_4;
    output akku_o_c_3;
    output akku_o_c_2;
    output akku_o_c_1;
    output \adrram[5] ;
    output \adrram[4] ;
    output \adrram[3] ;
    output \adrram[2] ;
    output \adrram[1] ;
    output n2313;
    input n2310;
    output we_N_63_enable_259;
    input n2314;
    output we_N_63_enable_315;
    input n2306;
    output we_N_63_enable_187;
    input reset_c;
    output we_N_63;
    output oe_N_57;
    output n2305;
    input GND_net;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/70735/desktop/cpu/cpu2system.vhd(9[13:16])
    wire we_N_63 /* synthesis is_clock=1, is_inv_clock=1, SET_AS_NETWORK=\CPU/we_N_63 */ ;   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(13[13:15])
    wire [5:0]adress_5__N_3;
    
    wire clk_c_enable_15;
    wire [8:0]akku_o_8__N_44;
    wire [5:0]pc;   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(23[15:17])
    
    wire clk_c_enable_7, n2304, n804;
    wire [5:0]pc_5__N_30_c;
    
    wire clk_c_enable_8;
    wire [8:0]akku_o_8__N_11;
    wire [2:0]states;   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(25[15:21])
    
    wire n2302, n2;
    wire [2:0]states_2__N_53;
    
    wire n2303, n2312;
    wire [7:0]akku_o_8__N_36;
    
    wire n1542, n1541, n1540, n1539, n1538;
    
    FD1S3AX adreg_i1 (.D(adress_5__N_3[0]), .CK(clk_c), .Q(\adrram[0] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=46, LSE_RLINE=46 */ ;   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(30[9] 71[16])
    defparam adreg_i1.GSR = "ENABLED";
    FD1P3AX akku_i1 (.D(akku_o_8__N_44[0]), .SP(clk_c_enable_15), .CK(clk_c), 
            .Q(akku_o_c_0)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=46, LSE_RLINE=46 */ ;   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(30[9] 71[16])
    defparam akku_i1.GSR = "ENABLED";
    FD1P3AX pc_i0_i0 (.D(pc_5__N_30[0]), .SP(clk_c_enable_7), .CK(clk_c), 
            .Q(pc[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=46, LSE_RLINE=46 */ ;   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(30[9] 71[16])
    defparam pc_i0_i0.GSR = "ENABLED";
    LUT4 i696_2_lut_3_lut_4_lut (.A(data[7]), .B(akku_o_c_8), .C(n2304), 
         .D(data[6]), .Z(n804)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;
    defparam i696_2_lut_3_lut_4_lut.init = 16'hf8f0;
    FD1P3AX pc_i0_i5 (.D(pc_5__N_30_c[5]), .SP(clk_c_enable_7), .CK(clk_c), 
            .Q(pc[5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=46, LSE_RLINE=46 */ ;   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(30[9] 71[16])
    defparam pc_i0_i5.GSR = "ENABLED";
    FD1P3AX pc_i0_i4 (.D(pc_5__N_30_c[4]), .SP(clk_c_enable_7), .CK(clk_c), 
            .Q(pc[4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=46, LSE_RLINE=46 */ ;   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(30[9] 71[16])
    defparam pc_i0_i4.GSR = "ENABLED";
    FD1P3AX pc_i0_i3 (.D(pc_5__N_30_c[3]), .SP(clk_c_enable_7), .CK(clk_c), 
            .Q(pc[3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=46, LSE_RLINE=46 */ ;   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(30[9] 71[16])
    defparam pc_i0_i3.GSR = "ENABLED";
    FD1P3AX pc_i0_i2 (.D(pc_5__N_30_c[2]), .SP(clk_c_enable_7), .CK(clk_c), 
            .Q(pc[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=46, LSE_RLINE=46 */ ;   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(30[9] 71[16])
    defparam pc_i0_i2.GSR = "ENABLED";
    FD1P3AX pc_i0_i1 (.D(pc_5__N_30_c[1]), .SP(clk_c_enable_7), .CK(clk_c), 
            .Q(pc[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=46, LSE_RLINE=46 */ ;   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(30[9] 71[16])
    defparam pc_i0_i1.GSR = "ENABLED";
    FD1P3AX akku_i9 (.D(akku_o_8__N_11[8]), .SP(clk_c_enable_8), .CK(clk_c), 
            .Q(akku_o_c_8)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=46, LSE_RLINE=46 */ ;   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(30[9] 71[16])
    defparam akku_i9.GSR = "ENABLED";
    FD1P3AX akku_i8 (.D(akku_o_8__N_44[7]), .SP(clk_c_enable_15), .CK(clk_c), 
            .Q(akku_o_c_7)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=46, LSE_RLINE=46 */ ;   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(30[9] 71[16])
    defparam akku_i8.GSR = "ENABLED";
    FD1P3AX akku_i7 (.D(akku_o_8__N_44[6]), .SP(clk_c_enable_15), .CK(clk_c), 
            .Q(akku_o_c_6)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=46, LSE_RLINE=46 */ ;   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(30[9] 71[16])
    defparam akku_i7.GSR = "ENABLED";
    FD1P3AX akku_i6 (.D(akku_o_8__N_44[5]), .SP(clk_c_enable_15), .CK(clk_c), 
            .Q(akku_o_c_5)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=46, LSE_RLINE=46 */ ;   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(30[9] 71[16])
    defparam akku_i6.GSR = "ENABLED";
    FD1P3AX akku_i5 (.D(akku_o_8__N_44[4]), .SP(clk_c_enable_15), .CK(clk_c), 
            .Q(akku_o_c_4)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=46, LSE_RLINE=46 */ ;   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(30[9] 71[16])
    defparam akku_i5.GSR = "ENABLED";
    FD1P3AX akku_i4 (.D(akku_o_8__N_44[3]), .SP(clk_c_enable_15), .CK(clk_c), 
            .Q(akku_o_c_3)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=46, LSE_RLINE=46 */ ;   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(30[9] 71[16])
    defparam akku_i4.GSR = "ENABLED";
    FD1P3AX akku_i3 (.D(akku_o_8__N_44[2]), .SP(clk_c_enable_15), .CK(clk_c), 
            .Q(akku_o_c_2)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=46, LSE_RLINE=46 */ ;   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(30[9] 71[16])
    defparam akku_i3.GSR = "ENABLED";
    FD1P3AX akku_i2 (.D(akku_o_8__N_44[1]), .SP(clk_c_enable_15), .CK(clk_c), 
            .Q(akku_o_c_1)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=46, LSE_RLINE=46 */ ;   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(30[9] 71[16])
    defparam akku_i2.GSR = "ENABLED";
    FD1S3AX adreg_i6 (.D(adress_5__N_3[5]), .CK(clk_c), .Q(\adrram[5] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=46, LSE_RLINE=46 */ ;   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(30[9] 71[16])
    defparam adreg_i6.GSR = "ENABLED";
    FD1S3AX adreg_i5 (.D(adress_5__N_3[4]), .CK(clk_c), .Q(\adrram[4] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=46, LSE_RLINE=46 */ ;   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(30[9] 71[16])
    defparam adreg_i5.GSR = "ENABLED";
    FD1S3AX adreg_i4 (.D(adress_5__N_3[3]), .CK(clk_c), .Q(\adrram[3] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=46, LSE_RLINE=46 */ ;   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(30[9] 71[16])
    defparam adreg_i4.GSR = "ENABLED";
    FD1S3AX adreg_i3 (.D(adress_5__N_3[2]), .CK(clk_c), .Q(\adrram[2] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=46, LSE_RLINE=46 */ ;   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(30[9] 71[16])
    defparam adreg_i3.GSR = "ENABLED";
    FD1S3AX adreg_i2 (.D(adress_5__N_3[1]), .CK(clk_c), .Q(\adrram[1] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=46, LSE_RLINE=46 */ ;   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(30[9] 71[16])
    defparam adreg_i2.GSR = "ENABLED";
    FD1S3IX states__i2 (.D(n2302), .CK(clk_c), .CD(n2304), .Q(states[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=46, LSE_RLINE=46 */ ;   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(30[9] 71[16])
    defparam states__i2.GSR = "ENABLED";
    FD1S3IX states__i1 (.D(n2), .CK(clk_c), .CD(n804), .Q(states[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=46, LSE_RLINE=46 */ ;   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(30[9] 71[16])
    defparam states__i1.GSR = "ENABLED";
    FD1S3IX states__i0 (.D(states_2__N_53[0]), .CK(clk_c), .CD(n2304), 
            .Q(states[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=46, LSE_RLINE=46 */ ;   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(30[9] 71[16])
    defparam states__i0.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_15_3_lut (.A(data[7]), .B(akku_o_c_8), .C(data[6]), 
         .Z(n2302)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_rep_15_3_lut.init = 16'h8080;
    LUT4 i1154_2_lut_3_lut (.A(data[7]), .B(akku_o_c_8), .C(data[6]), 
         .Z(states_2__N_53[0])) /* synthesis lut_function=(A (B+!(C))+!A !(C)) */ ;
    defparam i1154_2_lut_3_lut.init = 16'h8f8f;
    LUT4 i2278_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2313), .C(n2310), 
         .D(\adrram[5] ), .Z(we_N_63_enable_259)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // E:/Diamond/diamond/3.10_x64/ispfpga/vhdl_packages/numeric_std.vhd(1241[12:13])
    defparam i2278_2_lut_2_lut_3_lut_4_lut.init = 16'h0008;
    LUT4 i460_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2313), .C(\adrram[4] ), 
         .D(\adrram[3] ), .Z(pc_5__N_30_c[4])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // E:/Diamond/diamond/3.10_x64/ispfpga/vhdl_packages/numeric_std.vhd(1241[12:13])
    defparam i460_2_lut_3_lut_4_lut.init = 16'h78f0;
    LUT4 i2240_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2313), .C(n2314), 
         .D(\adrram[5] ), .Z(we_N_63_enable_315)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // E:/Diamond/diamond/3.10_x64/ispfpga/vhdl_packages/numeric_std.vhd(1241[12:13])
    defparam i2240_2_lut_2_lut_3_lut_4_lut.init = 16'h0008;
    LUT4 i2342_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2313), .C(n2306), 
         .D(\adrram[5] ), .Z(we_N_63_enable_187)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // E:/Diamond/diamond/3.10_x64/ispfpga/vhdl_packages/numeric_std.vhd(1241[12:13])
    defparam i2342_2_lut_2_lut_3_lut_4_lut.init = 16'h0080;
    LUT4 i467_3_lut_4_lut (.A(\adrram[3] ), .B(n2303), .C(\adrram[4] ), 
         .D(\adrram[5] ), .Z(pc_5__N_30_c[5])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // E:/Diamond/diamond/3.10_x64/ispfpga/vhdl_packages/numeric_std.vhd(1241[12:13])
    defparam i467_3_lut_4_lut.init = 16'h7f80;
    LUT4 pc_5__I_0_85_i3_3_lut_4_lut (.A(states[0]), .B(n2312), .C(pc[2]), 
         .D(data[2]), .Z(adress_5__N_3[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(76[33:48])
    defparam pc_5__I_0_85_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 pc_5__I_0_85_i1_3_lut_4_lut (.A(states[0]), .B(n2312), .C(pc[0]), 
         .D(data[0]), .Z(adress_5__N_3[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(76[33:48])
    defparam pc_5__I_0_85_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 pc_5__I_0_85_i6_3_lut_4_lut (.A(states[0]), .B(n2312), .C(pc[5]), 
         .D(data[5]), .Z(adress_5__N_3[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(76[33:48])
    defparam pc_5__I_0_85_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 pc_5__I_0_85_i5_3_lut_4_lut (.A(states[0]), .B(n2312), .C(pc[4]), 
         .D(data[4]), .Z(adress_5__N_3[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(76[33:48])
    defparam pc_5__I_0_85_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 pc_5__I_0_85_i4_3_lut_4_lut (.A(states[0]), .B(n2312), .C(pc[3]), 
         .D(data[3]), .Z(adress_5__N_3[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(76[33:48])
    defparam pc_5__I_0_85_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 pc_5__I_0_85_i2_3_lut_4_lut (.A(states[0]), .B(n2312), .C(pc[1]), 
         .D(data[1]), .Z(adress_5__N_3[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(76[33:48])
    defparam pc_5__I_0_85_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i439_2_lut (.A(\adrram[1] ), .B(\adrram[0] ), .Z(pc_5__N_30_c[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // E:/Diamond/diamond/3.10_x64/ispfpga/vhdl_packages/numeric_std.vhd(1241[12:13])
    defparam i439_2_lut.init = 16'h6666;
    LUT4 i1159_2_lut (.A(akku_o_8__N_44[8]), .B(states[2]), .Z(akku_o_8__N_11[8])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(47[13] 54[22])
    defparam i1159_2_lut.init = 16'h2222;
    LUT4 i482_1_lut (.A(data[7]), .Z(n2)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(59[20:43])
    defparam i482_1_lut.init = 16'h5555;
    LUT4 i2252_2_lut (.A(akku_o_c_6), .B(data[6]), .Z(akku_o_8__N_36[6])) /* synthesis lut_function=(!(A+(B))) */ ;   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(50[60:94])
    defparam i2252_2_lut.init = 16'h1111;
    LUT4 i2249_2_lut (.A(akku_o_c_7), .B(data[7]), .Z(akku_o_8__N_36[7])) /* synthesis lut_function=(!(A+(B))) */ ;   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(50[60:94])
    defparam i2249_2_lut.init = 16'h1111;
    LUT4 i2258_2_lut (.A(akku_o_c_4), .B(data[4]), .Z(akku_o_8__N_36[4])) /* synthesis lut_function=(!(A+(B))) */ ;   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(50[60:94])
    defparam i2258_2_lut.init = 16'h1111;
    LUT4 i2255_2_lut (.A(akku_o_c_5), .B(data[5]), .Z(akku_o_8__N_36[5])) /* synthesis lut_function=(!(A+(B))) */ ;   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(50[60:94])
    defparam i2255_2_lut.init = 16'h1111;
    LUT4 i2264_2_lut (.A(akku_o_c_2), .B(data[2]), .Z(akku_o_8__N_36[2])) /* synthesis lut_function=(!(A+(B))) */ ;   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(50[60:94])
    defparam i2264_2_lut.init = 16'h1111;
    LUT4 i2261_2_lut (.A(akku_o_c_3), .B(data[3]), .Z(akku_o_8__N_36[3])) /* synthesis lut_function=(!(A+(B))) */ ;   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(50[60:94])
    defparam i2261_2_lut.init = 16'h1111;
    LUT4 i2270_2_lut (.A(akku_o_c_0), .B(data[0]), .Z(akku_o_8__N_36[0])) /* synthesis lut_function=(!(A+(B))) */ ;   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(50[60:94])
    defparam i2270_2_lut.init = 16'h1111;
    LUT4 i2267_2_lut (.A(akku_o_c_1), .B(data[1]), .Z(akku_o_8__N_36[1])) /* synthesis lut_function=(!(A+(B))) */ ;   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(50[60:94])
    defparam i2267_2_lut.init = 16'h1111;
    LUT4 i703_2_lut_rep_24 (.A(states[1]), .B(states[2]), .Z(clk_c_enable_15)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(47[13] 54[22])
    defparam i703_2_lut_rep_24.init = 16'h2222;
    LUT4 i13_4_lut_3_lut (.A(states[1]), .B(states[2]), .C(states[0]), 
         .Z(clk_c_enable_8)) /* synthesis lut_function=(!(A (B+(C))+!A !(B (C)))) */ ;   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(47[13] 54[22])
    defparam i13_4_lut_3_lut.init = 16'h4242;
    LUT4 i2203_2_lut_2_lut_3_lut_4_lut (.A(reset_c), .B(clk_c), .C(n2312), 
         .D(states[0]), .Z(we_N_63)) /* synthesis lut_function=((B+(C+!(D)))+!A) */ ;   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(82[21:60])
    defparam i2203_2_lut_2_lut_3_lut_4_lut.init = 16'hfdff;
    LUT4 i1_3_lut_4_lut (.A(reset_c), .B(clk_c), .C(states[1]), .D(states[0]), 
         .Z(oe_N_57)) /* synthesis lut_function=(!((B+!(C+!(D)))+!A)) */ ;   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(82[21:60])
    defparam i1_3_lut_4_lut.init = 16'h2022;
    LUT4 i1_2_lut_rep_25 (.A(states[1]), .B(states[2]), .Z(n2312)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(76[33:48])
    defparam i1_2_lut_rep_25.init = 16'heeee;
    LUT4 i1_2_lut_rep_17_3_lut (.A(states[1]), .B(states[2]), .C(states[0]), 
         .Z(n2304)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(76[33:48])
    defparam i1_2_lut_rep_17_3_lut.init = 16'hfefe;
    LUT4 i834_1_lut_2_lut_3_lut (.A(states[1]), .B(states[2]), .C(states[0]), 
         .Z(clk_c_enable_7)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(76[33:48])
    defparam i834_1_lut_2_lut_3_lut.init = 16'h0101;
    LUT4 i1_2_lut_rep_18_3_lut (.A(states[1]), .B(states[2]), .C(states[0]), 
         .Z(n2305)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(76[33:48])
    defparam i1_2_lut_rep_18_3_lut.init = 16'hefef;
    LUT4 i441_2_lut_rep_26 (.A(\adrram[1] ), .B(\adrram[0] ), .Z(n2313)) /* synthesis lut_function=(A (B)) */ ;   // E:/Diamond/diamond/3.10_x64/ispfpga/vhdl_packages/numeric_std.vhd(1241[12:13])
    defparam i441_2_lut_rep_26.init = 16'h8888;
    LUT4 i448_2_lut_rep_16_3_lut (.A(\adrram[1] ), .B(\adrram[0] ), .C(\adrram[2] ), 
         .Z(n2303)) /* synthesis lut_function=(A (B (C))) */ ;   // E:/Diamond/diamond/3.10_x64/ispfpga/vhdl_packages/numeric_std.vhd(1241[12:13])
    defparam i448_2_lut_rep_16_3_lut.init = 16'h8080;
    LUT4 i446_2_lut_3_lut (.A(\adrram[1] ), .B(\adrram[0] ), .C(\adrram[2] ), 
         .Z(pc_5__N_30_c[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // E:/Diamond/diamond/3.10_x64/ispfpga/vhdl_packages/numeric_std.vhd(1241[12:13])
    defparam i446_2_lut_3_lut.init = 16'h7878;
    LUT4 i453_2_lut_3_lut_4_lut (.A(\adrram[1] ), .B(\adrram[0] ), .C(\adrram[3] ), 
         .D(\adrram[2] ), .Z(pc_5__N_30_c[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // E:/Diamond/diamond/3.10_x64/ispfpga/vhdl_packages/numeric_std.vhd(1241[12:13])
    defparam i453_2_lut_3_lut_4_lut.init = 16'h78f0;
    CCU2D add_91_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n1542), 
          .S0(akku_o_8__N_44[8]));   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(48[39:69])
    defparam add_91_cout.INIT0 = 16'h0000;
    defparam add_91_cout.INIT1 = 16'h0000;
    defparam add_91_cout.INJECT1_0 = "NO";
    defparam add_91_cout.INJECT1_1 = "NO";
    CCU2D add_91_9 (.A0(data[6]), .B0(states[0]), .C0(akku_o_8__N_36[6]), 
          .D0(akku_o_c_6), .A1(data[7]), .B1(states[0]), .C1(akku_o_8__N_36[7]), 
          .D1(akku_o_c_7), .CIN(n1541), .COUT(n1542), .S0(akku_o_8__N_44[6]), 
          .S1(akku_o_8__N_44[7]));   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(48[39:69])
    defparam add_91_9.INIT0 = 16'hd1e2;
    defparam add_91_9.INIT1 = 16'hd1e2;
    defparam add_91_9.INJECT1_0 = "NO";
    defparam add_91_9.INJECT1_1 = "NO";
    CCU2D add_91_7 (.A0(data[4]), .B0(states[0]), .C0(akku_o_8__N_36[4]), 
          .D0(akku_o_c_4), .A1(data[5]), .B1(states[0]), .C1(akku_o_8__N_36[5]), 
          .D1(akku_o_c_5), .CIN(n1540), .COUT(n1541), .S0(akku_o_8__N_44[4]), 
          .S1(akku_o_8__N_44[5]));   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(48[39:69])
    defparam add_91_7.INIT0 = 16'hd1e2;
    defparam add_91_7.INIT1 = 16'hd1e2;
    defparam add_91_7.INJECT1_0 = "NO";
    defparam add_91_7.INJECT1_1 = "NO";
    CCU2D add_91_5 (.A0(data[2]), .B0(states[0]), .C0(akku_o_8__N_36[2]), 
          .D0(akku_o_c_2), .A1(data[3]), .B1(states[0]), .C1(akku_o_8__N_36[3]), 
          .D1(akku_o_c_3), .CIN(n1539), .COUT(n1540), .S0(akku_o_8__N_44[2]), 
          .S1(akku_o_8__N_44[3]));   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(48[39:69])
    defparam add_91_5.INIT0 = 16'hd1e2;
    defparam add_91_5.INIT1 = 16'hd1e2;
    defparam add_91_5.INJECT1_0 = "NO";
    defparam add_91_5.INJECT1_1 = "NO";
    CCU2D add_91_3 (.A0(data[0]), .B0(states[0]), .C0(akku_o_8__N_36[0]), 
          .D0(akku_o_c_0), .A1(data[1]), .B1(states[0]), .C1(akku_o_8__N_36[1]), 
          .D1(akku_o_c_1), .CIN(n1538), .COUT(n1539), .S0(akku_o_8__N_44[0]), 
          .S1(akku_o_8__N_44[1]));   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(48[39:69])
    defparam add_91_3.INIT0 = 16'hd1e2;
    defparam add_91_3.INIT1 = 16'hd1e2;
    defparam add_91_3.INJECT1_0 = "NO";
    defparam add_91_3.INJECT1_1 = "NO";
    CCU2D add_91_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(states[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n1538));   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(48[39:69])
    defparam add_91_1.INIT0 = 16'hF000;
    defparam add_91_1.INIT1 = 16'h0fff;
    defparam add_91_1.INJECT1_0 = "NO";
    defparam add_91_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module TSALL
// module not written out since it is a black-box. 
//

//
// Verilog Description of module sram64kx8
//

module sram64kx8 (we_N_63, data, we_N_63_enable_315, we_N_63_enable_259, 
            we_N_63_enable_187, akku_o_c_0, oe_N_57, n2305, akku_o_c_5, 
            \adrram[0] , \adrram[2] , n2314, \adrram[5] , \adrram[3] , 
            \adrram[1] , n2306, n2310, akku_o_c_4, akku_o_c_3, n2313, 
            \pc_5__N_30[0] , \adrram[4] , akku_o_c_6, akku_o_c_2, akku_o_c_1, 
            akku_o_c_7);
    input we_N_63;
    output [7:0]data;
    input we_N_63_enable_315;
    input we_N_63_enable_259;
    input we_N_63_enable_187;
    input akku_o_c_0;
    input oe_N_57;
    input n2305;
    input akku_o_c_5;
    input \adrram[0] ;
    input \adrram[2] ;
    output n2314;
    input \adrram[5] ;
    input \adrram[3] ;
    input \adrram[1] ;
    output n2306;
    output n2310;
    input akku_o_c_4;
    input akku_o_c_3;
    input n2313;
    output \pc_5__N_30[0] ;
    input \adrram[4] ;
    input akku_o_c_6;
    input akku_o_c_2;
    input akku_o_c_1;
    input akku_o_c_7;
    
    wire we_N_63 /* synthesis is_clock=1, is_inv_clock=1, SET_AS_NETWORK=\CPU/we_N_63 */ ;   // c:/users/70735/desktop/cpu/tb02cpu2.vhd(13[13:15])
    wire [7:0]\mem[2] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_481;
    wire [7:0]\mem[1] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_452;
    wire [7:0]\mem[43] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_219;
    wire [7:0]\mem[50] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_512;
    wire [7:0]\mem[42] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_137;
    wire [7:0]\mem[3] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_416;
    wire [7:0]\mem[41] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_136;
    wire [7:0]\mem[40] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_135;
    wire [7:0]\mem[39] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_134;
    wire [7:0]\mem[49] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_144;
    wire [7:0]\mem[38] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_133;
    wire [7:0]\mem[37] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_132;
    wire [7:0]\mem[36] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_131;
    wire [7:0]\mem[35] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_130;
    wire [7:0]\mem[48] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_143;
    wire [7:0]\mem[34] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_129;
    wire [7:0]\mem[33] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_160;
    wire [7:0]\mem[4] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_407;
    wire [7:0]\mem[5] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_395;
    wire [7:0]\mem[6] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_386;
    wire [7:0]\mem[7] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_377;
    wire [7:0]\mem[8] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_368;
    wire [7:0]\mem[9] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_359;
    wire [7:0]\mem[10] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_351;
    wire [7:0]\mem[11] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_343;
    wire [7:0]\mem[12] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_336;
    wire [7:0]\mem[13] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_329;
    wire [7:0]\mem[14] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_322;
    wire [7:0]\mem[15] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    wire [7:0]\mem[16] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_308;
    wire [7:0]\mem[17] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_301;
    wire [7:0]\mem[18] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_294;
    wire [7:0]\mem[19] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_287;
    wire [7:0]\mem[20] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_280;
    wire [7:0]\mem[21] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_273;
    wire [7:0]\mem[22] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_266;
    wire [7:0]\mem[23] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    wire [7:0]\mem[24] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_252;
    wire [7:0]\mem[25] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_245;
    wire [7:0]\mem[26] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_238;
    wire [7:0]\mem[27] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_231;
    wire [7:0]\mem[28] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_224;
    wire [7:0]\mem[29] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_216;
    wire [7:0]\mem[30] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_201;
    wire [7:0]\mem[31] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    wire [7:0]\mem[32] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_173;
    wire [7:0]\mem[44] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_213;
    wire [7:0]\mem[45] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_202;
    wire [7:0]\mem[46] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_188;
    wire [7:0]\mem[47] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_174;
    wire [7:0]\mem[51] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_511;
    wire [7:0]\mem[52] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_504;
    wire [7:0]\mem[53] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_497;
    wire [7:0]\mem[54] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_490;
    wire [7:0]\mem[55] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_483;
    wire [7:0]\mem[56] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_474;
    wire [7:0]\mem[57] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_465;
    wire [7:0]\mem[58] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_455;
    wire [7:0]\mem[59] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_446;
    wire [7:0]\mem[60] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_437;
    wire [7:0]\mem[61] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_428;
    wire [7:0]\mem[62] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_420;
    wire [7:0]\mem[63] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_405;
    wire [7:0]\mem[0] ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(50[12:15])
    
    wire we_N_63_enable_379;
    wire [7:0]data_7__N_66;
    
    wire n1904, n1903, n2005, n2004, n1902, n1901, n2003, n2002, 
        n2001, n2000, n1999, n1998, n1602, n1601, n1997, n1996, 
        n1995, n1994, n1600, n1599, n1598, n1597, n1596, n1595, 
        n1699, n1698, n1594, n1593, n1697, n1696, n1695, n1694, 
        n1693, n1692, n1691, n1690, n1822, n2065, n1947, n2067, 
        n2064, n1946, n1936, n2066, n2063, n2059, n1821, n2062, 
        n2058, n1935, n1820, n1934, n1753, n1716, n1792, n1945, 
        n1752, n2307, n2030, n1791, n1944, n1933, n1715, n1635, 
        n2029, n1932, n1751, n1634, n2061, n1943, n1750, n1916, 
        n2028, n2060, n1942, n1761, n1915, n1633, n1908, n1689, 
        n2027, n1790, n1838, n1869, n1807, n1900, n1789, n1776, 
        n1931, n1745, n1962, n1714, n1993, n1819, n1683, n2024, 
        n1652, n2055, n1621, n2086, n1677, n1678, n1681, n1818, 
        n1679, n1680, n1682, n1615, n1616, n1619, n1741, n1742, 
        n1744, n1739, n1740, n1743, n1863, n1864, n1867, n1941, 
        n1865, n1866, n1868, n1987, n1988, n1991, n1989, n1990, 
        n1992, n2049, n2050, n2053, n1760, n2051, n2052, n2054, 
        n2080, n2081, n2084, n2082, n2083, n2085, n1894, n1895, 
        n1898, n1788, n1896, n1897, n1899, n1646, n1647, n1650, 
        n1648, n1649, n1651, n1617, n1618, n1620, n1817, n1708, 
        n1709, n1712, n1787, n2068, n2069, n2078, n1636, n1637, 
        n1645, n1940, n1816, n1786, n1749, n1785, n1815, n1814, 
        n1939, n1759, n1784, n1813, n1783, n1938, n1758, n1748, 
        n1812, n1782, n1781, n1811, n1810, n2057, n1963, n1964, 
        n1979, n1757, n1747, n1604, n1632, n1780, n1809, n1779, 
        n2056, n1756, n1746, n1603, n1907, n1808, n1778, n1912, 
        n1777, n2026, n2025, n1937, n1755, n1718, n1914, n1911, 
        n1688, n1847, n1848, n1977, n1978, n1849, n1850, n1851, 
        n1852, n1853, n1854, n1729, n1730, n1727, n1728, n1725, 
        n1726, n1723, n1724, n1721, n1722, n1719, n1720, n1591, 
        n1592, n1754, n1717, n2007, n2009, n2008, n1631, n1630, 
        n1687, n1686, n1685, n1684, n1885, n1884, n1883, n1882, 
        n1881, n1880, n1910, n1909, n2006, n1629, n1628, n1625, 
        n1624, n1623, n1913, n1627, n1622, n1626, n1906, n1905, 
        n1879, n1878, n1877, n1876, n1875, n1874, n1873, n1872, 
        n1871, n1870, n1846, n2031, n2032, n2044, n1845, n1976, 
        n1975, n1844, n1843, n1842, n1841, n1974, n1973, n2040, 
        n2039, n1840, n1839, n1972, n1971, n1970, n1969, n2038, 
        n2037, n1968, n1967, n1668, n1667, n1666, n1665, n1966, 
        n1965, n2036, n2035, n2071, n2070, n1606, n1605, n1664, 
        n1663, n1662, n1661, n1660, n1659, n1658, n1657, n1656, 
        n1655, n1654, n1653, n2315, n2309, n2308, n2033, n2034, 
        n2045, n1710, n1711, n1713, n1925, n1926, n1929, n1927, 
        n1928, n1930, n2018, n2019, n2022, n2020, n2021, n2023, 
        n1770, n1771, n1774, n1772, n1773, n1775, n1801, n1802, 
        n1805, n1803, n1804, n1806, n1956, n1957, n1960, n1958, 
        n1959, n1961, n1832, n1833, n1836, n1834, n1835, n1837, 
        n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, 
        n1611, n1612, n2072, n2073, n1613, n1614, n2041, n2042, 
        n1980, n1855, n1856, n2074, n2075, n2043, n1981, n1982, 
        n1857, n1858, n1859, n1860, n1737, n1738, n1735, n1736, 
        n1983, n1984, n1861, n1862, n1733, n1734, n1731, n1732, 
        n2046, n1985, n1986, n2076, n2077, n2047, n2048, n2079, 
        n1638, n1639, n1640, n1641, n1642, n1643, n1886, n1887, 
        n1888, n1889, n1890, n1891, n1892, n1893, n1644, n1700, 
        n1701, n2010, n2011, n1702, n1703, n1704, n1705, n1917, 
        n1918, n1706, n1707, n2012, n2013, n1919, n1920, n1921, 
        n1922, n2014, n2015, n1923, n1924, n2016, n2017, n1762, 
        n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1948, 
        n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1793, 
        n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1609, 
        n1610, n1824, n1825, n1826, n1827, n1828, n1829, n1830, 
        n1831, n1607, n1608, n1823;
    
    FD1P3AY mem_2__i0_i0 (.D(data[0]), .SP(we_N_63_enable_481), .CK(we_N_63), 
            .Q(\mem[2] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_2__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_1__i0_i0 (.D(data[0]), .SP(we_N_63_enable_452), .CK(we_N_63), 
            .Q(\mem[1] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_1__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_43__i0_i5 (.D(data[5]), .SP(we_N_63_enable_219), .CK(we_N_63), 
            .Q(\mem[43] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_43__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_43__i0_i4 (.D(data[4]), .SP(we_N_63_enable_219), .CK(we_N_63), 
            .Q(\mem[43] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_43__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_43__i0_i3 (.D(data[3]), .SP(we_N_63_enable_219), .CK(we_N_63), 
            .Q(\mem[43] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_43__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_50__i0_i6 (.D(data[6]), .SP(we_N_63_enable_512), .CK(we_N_63), 
            .Q(\mem[50] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_50__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_50__i0_i5 (.D(data[5]), .SP(we_N_63_enable_512), .CK(we_N_63), 
            .Q(\mem[50] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_50__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_50__i0_i4 (.D(data[4]), .SP(we_N_63_enable_512), .CK(we_N_63), 
            .Q(\mem[50] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_50__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_43__i0_i2 (.D(data[2]), .SP(we_N_63_enable_219), .CK(we_N_63), 
            .Q(\mem[43] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_43__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_50__i0_i3 (.D(data[3]), .SP(we_N_63_enable_512), .CK(we_N_63), 
            .Q(\mem[50] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_50__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_43__i0_i1 (.D(data[1]), .SP(we_N_63_enable_219), .CK(we_N_63), 
            .Q(\mem[43] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_43__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_50__i0_i2 (.D(data[2]), .SP(we_N_63_enable_512), .CK(we_N_63), 
            .Q(\mem[50] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_50__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_42__i0_i7 (.D(data[7]), .SP(we_N_63_enable_137), .CK(we_N_63), 
            .Q(\mem[42] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_42__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_42__i0_i6 (.D(data[6]), .SP(we_N_63_enable_137), .CK(we_N_63), 
            .Q(\mem[42] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_42__i0_i6.GSR = "ENABLED";
    FD1P3AY mem_3__i0_i0 (.D(data[0]), .SP(we_N_63_enable_416), .CK(we_N_63), 
            .Q(\mem[3] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_3__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_42__i0_i5 (.D(data[5]), .SP(we_N_63_enable_137), .CK(we_N_63), 
            .Q(\mem[42] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_42__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_42__i0_i4 (.D(data[4]), .SP(we_N_63_enable_137), .CK(we_N_63), 
            .Q(\mem[42] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_42__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_42__i0_i3 (.D(data[3]), .SP(we_N_63_enable_137), .CK(we_N_63), 
            .Q(\mem[42] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_42__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_42__i0_i2 (.D(data[2]), .SP(we_N_63_enable_137), .CK(we_N_63), 
            .Q(\mem[42] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_42__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_42__i0_i1 (.D(data[1]), .SP(we_N_63_enable_137), .CK(we_N_63), 
            .Q(\mem[42] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_42__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_41__i0_i7 (.D(data[7]), .SP(we_N_63_enable_136), .CK(we_N_63), 
            .Q(\mem[41] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_41__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_41__i0_i6 (.D(data[6]), .SP(we_N_63_enable_136), .CK(we_N_63), 
            .Q(\mem[41] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_41__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_41__i0_i5 (.D(data[5]), .SP(we_N_63_enable_136), .CK(we_N_63), 
            .Q(\mem[41] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_41__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_41__i0_i4 (.D(data[4]), .SP(we_N_63_enable_136), .CK(we_N_63), 
            .Q(\mem[41] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_41__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_41__i0_i3 (.D(data[3]), .SP(we_N_63_enable_136), .CK(we_N_63), 
            .Q(\mem[41] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_41__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_41__i0_i2 (.D(data[2]), .SP(we_N_63_enable_136), .CK(we_N_63), 
            .Q(\mem[41] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_41__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_41__i0_i1 (.D(data[1]), .SP(we_N_63_enable_136), .CK(we_N_63), 
            .Q(\mem[41] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_41__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_40__i0_i7 (.D(data[7]), .SP(we_N_63_enable_135), .CK(we_N_63), 
            .Q(\mem[40] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_40__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_40__i0_i6 (.D(data[6]), .SP(we_N_63_enable_135), .CK(we_N_63), 
            .Q(\mem[40] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_40__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_40__i0_i5 (.D(data[5]), .SP(we_N_63_enable_135), .CK(we_N_63), 
            .Q(\mem[40] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_40__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_40__i0_i4 (.D(data[4]), .SP(we_N_63_enable_135), .CK(we_N_63), 
            .Q(\mem[40] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_40__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_40__i0_i3 (.D(data[3]), .SP(we_N_63_enable_135), .CK(we_N_63), 
            .Q(\mem[40] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_40__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_40__i0_i2 (.D(data[2]), .SP(we_N_63_enable_135), .CK(we_N_63), 
            .Q(\mem[40] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_40__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_50__i0_i1 (.D(data[1]), .SP(we_N_63_enable_512), .CK(we_N_63), 
            .Q(\mem[50] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_50__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_40__i0_i1 (.D(data[1]), .SP(we_N_63_enable_135), .CK(we_N_63), 
            .Q(\mem[40] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_40__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_39__i0_i7 (.D(data[7]), .SP(we_N_63_enable_134), .CK(we_N_63), 
            .Q(\mem[39] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_39__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_49__i0_i7 (.D(data[7]), .SP(we_N_63_enable_144), .CK(we_N_63), 
            .Q(\mem[49] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_49__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_39__i0_i6 (.D(data[6]), .SP(we_N_63_enable_134), .CK(we_N_63), 
            .Q(\mem[39] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_39__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_43__i0_i6 (.D(data[6]), .SP(we_N_63_enable_219), .CK(we_N_63), 
            .Q(\mem[43] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_43__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_39__i0_i5 (.D(data[5]), .SP(we_N_63_enable_134), .CK(we_N_63), 
            .Q(\mem[39] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_39__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_39__i0_i4 (.D(data[4]), .SP(we_N_63_enable_134), .CK(we_N_63), 
            .Q(\mem[39] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_39__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_39__i0_i3 (.D(data[3]), .SP(we_N_63_enable_134), .CK(we_N_63), 
            .Q(\mem[39] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_39__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_39__i0_i2 (.D(data[2]), .SP(we_N_63_enable_134), .CK(we_N_63), 
            .Q(\mem[39] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_39__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_49__i0_i6 (.D(data[6]), .SP(we_N_63_enable_144), .CK(we_N_63), 
            .Q(\mem[49] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_49__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_39__i0_i1 (.D(data[1]), .SP(we_N_63_enable_134), .CK(we_N_63), 
            .Q(\mem[39] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_39__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_38__i0_i7 (.D(data[7]), .SP(we_N_63_enable_133), .CK(we_N_63), 
            .Q(\mem[38] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_38__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_38__i0_i6 (.D(data[6]), .SP(we_N_63_enable_133), .CK(we_N_63), 
            .Q(\mem[38] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_38__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_38__i0_i5 (.D(data[5]), .SP(we_N_63_enable_133), .CK(we_N_63), 
            .Q(\mem[38] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_38__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_38__i0_i4 (.D(data[4]), .SP(we_N_63_enable_133), .CK(we_N_63), 
            .Q(\mem[38] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_38__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_38__i0_i3 (.D(data[3]), .SP(we_N_63_enable_133), .CK(we_N_63), 
            .Q(\mem[38] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_38__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_38__i0_i2 (.D(data[2]), .SP(we_N_63_enable_133), .CK(we_N_63), 
            .Q(\mem[38] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_38__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_49__i0_i5 (.D(data[5]), .SP(we_N_63_enable_144), .CK(we_N_63), 
            .Q(\mem[49] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_49__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_38__i0_i1 (.D(data[1]), .SP(we_N_63_enable_133), .CK(we_N_63), 
            .Q(\mem[38] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_38__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_37__i0_i7 (.D(data[7]), .SP(we_N_63_enable_132), .CK(we_N_63), 
            .Q(\mem[37] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_37__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_37__i0_i6 (.D(data[6]), .SP(we_N_63_enable_132), .CK(we_N_63), 
            .Q(\mem[37] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_37__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_37__i0_i5 (.D(data[5]), .SP(we_N_63_enable_132), .CK(we_N_63), 
            .Q(\mem[37] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_37__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_37__i0_i4 (.D(data[4]), .SP(we_N_63_enable_132), .CK(we_N_63), 
            .Q(\mem[37] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_37__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_37__i0_i3 (.D(data[3]), .SP(we_N_63_enable_132), .CK(we_N_63), 
            .Q(\mem[37] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_37__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_37__i0_i2 (.D(data[2]), .SP(we_N_63_enable_132), .CK(we_N_63), 
            .Q(\mem[37] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_37__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_49__i0_i4 (.D(data[4]), .SP(we_N_63_enable_144), .CK(we_N_63), 
            .Q(\mem[49] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_49__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_37__i0_i1 (.D(data[1]), .SP(we_N_63_enable_132), .CK(we_N_63), 
            .Q(\mem[37] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_37__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_36__i0_i7 (.D(data[7]), .SP(we_N_63_enable_131), .CK(we_N_63), 
            .Q(\mem[36] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_36__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_36__i0_i6 (.D(data[6]), .SP(we_N_63_enable_131), .CK(we_N_63), 
            .Q(\mem[36] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_36__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_36__i0_i5 (.D(data[5]), .SP(we_N_63_enable_131), .CK(we_N_63), 
            .Q(\mem[36] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_36__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_36__i0_i4 (.D(data[4]), .SP(we_N_63_enable_131), .CK(we_N_63), 
            .Q(\mem[36] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_36__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_36__i0_i3 (.D(data[3]), .SP(we_N_63_enable_131), .CK(we_N_63), 
            .Q(\mem[36] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_36__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_36__i0_i2 (.D(data[2]), .SP(we_N_63_enable_131), .CK(we_N_63), 
            .Q(\mem[36] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_36__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_36__i0_i1 (.D(data[1]), .SP(we_N_63_enable_131), .CK(we_N_63), 
            .Q(\mem[36] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_36__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_35__i0_i7 (.D(data[7]), .SP(we_N_63_enable_130), .CK(we_N_63), 
            .Q(\mem[35] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_35__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_49__i0_i3 (.D(data[3]), .SP(we_N_63_enable_144), .CK(we_N_63), 
            .Q(\mem[49] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_49__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_49__i0_i2 (.D(data[2]), .SP(we_N_63_enable_144), .CK(we_N_63), 
            .Q(\mem[49] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_49__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_49__i0_i1 (.D(data[1]), .SP(we_N_63_enable_144), .CK(we_N_63), 
            .Q(\mem[49] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_49__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_35__i0_i6 (.D(data[6]), .SP(we_N_63_enable_130), .CK(we_N_63), 
            .Q(\mem[35] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_35__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_35__i0_i5 (.D(data[5]), .SP(we_N_63_enable_130), .CK(we_N_63), 
            .Q(\mem[35] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_35__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_35__i0_i4 (.D(data[4]), .SP(we_N_63_enable_130), .CK(we_N_63), 
            .Q(\mem[35] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_35__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_35__i0_i3 (.D(data[3]), .SP(we_N_63_enable_130), .CK(we_N_63), 
            .Q(\mem[35] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_35__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_35__i0_i2 (.D(data[2]), .SP(we_N_63_enable_130), .CK(we_N_63), 
            .Q(\mem[35] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_35__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_48__i0_i7 (.D(data[7]), .SP(we_N_63_enable_143), .CK(we_N_63), 
            .Q(\mem[48] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_48__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_48__i0_i6 (.D(data[6]), .SP(we_N_63_enable_143), .CK(we_N_63), 
            .Q(\mem[48] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_48__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_48__i0_i5 (.D(data[5]), .SP(we_N_63_enable_143), .CK(we_N_63), 
            .Q(\mem[48] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_48__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_35__i0_i1 (.D(data[1]), .SP(we_N_63_enable_130), .CK(we_N_63), 
            .Q(\mem[35] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_35__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_34__i0_i7 (.D(data[7]), .SP(we_N_63_enable_129), .CK(we_N_63), 
            .Q(\mem[34] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_34__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_34__i0_i6 (.D(data[6]), .SP(we_N_63_enable_129), .CK(we_N_63), 
            .Q(\mem[34] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_34__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_34__i0_i5 (.D(data[5]), .SP(we_N_63_enable_129), .CK(we_N_63), 
            .Q(\mem[34] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_34__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_34__i0_i4 (.D(data[4]), .SP(we_N_63_enable_129), .CK(we_N_63), 
            .Q(\mem[34] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_34__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_48__i0_i4 (.D(data[4]), .SP(we_N_63_enable_143), .CK(we_N_63), 
            .Q(\mem[48] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_48__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_48__i0_i3 (.D(data[3]), .SP(we_N_63_enable_143), .CK(we_N_63), 
            .Q(\mem[48] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_48__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_34__i0_i3 (.D(data[3]), .SP(we_N_63_enable_129), .CK(we_N_63), 
            .Q(\mem[34] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_34__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_34__i0_i2 (.D(data[2]), .SP(we_N_63_enable_129), .CK(we_N_63), 
            .Q(\mem[34] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_34__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_34__i0_i1 (.D(data[1]), .SP(we_N_63_enable_129), .CK(we_N_63), 
            .Q(\mem[34] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_34__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_33__i0_i7 (.D(data[7]), .SP(we_N_63_enable_160), .CK(we_N_63), 
            .Q(\mem[33] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_33__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_33__i0_i6 (.D(data[6]), .SP(we_N_63_enable_160), .CK(we_N_63), 
            .Q(\mem[33] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_33__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_33__i0_i5 (.D(data[5]), .SP(we_N_63_enable_160), .CK(we_N_63), 
            .Q(\mem[33] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_33__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_48__i0_i2 (.D(data[2]), .SP(we_N_63_enable_143), .CK(we_N_63), 
            .Q(\mem[48] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_48__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_48__i0_i1 (.D(data[1]), .SP(we_N_63_enable_143), .CK(we_N_63), 
            .Q(\mem[48] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_48__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_33__i0_i4 (.D(data[4]), .SP(we_N_63_enable_160), .CK(we_N_63), 
            .Q(\mem[33] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_33__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_33__i0_i3 (.D(data[3]), .SP(we_N_63_enable_160), .CK(we_N_63), 
            .Q(\mem[33] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_33__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_33__i0_i2 (.D(data[2]), .SP(we_N_63_enable_160), .CK(we_N_63), 
            .Q(\mem[33] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_33__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_4__i0_i0 (.D(data[0]), .SP(we_N_63_enable_407), .CK(we_N_63), 
            .Q(\mem[4] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_4__i0_i0.GSR = "ENABLED";
    FD1P3AY mem_5__i0_i0 (.D(data[0]), .SP(we_N_63_enable_395), .CK(we_N_63), 
            .Q(\mem[5] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_5__i0_i0.GSR = "ENABLED";
    FD1P3AY mem_6__i0_i0 (.D(data[0]), .SP(we_N_63_enable_386), .CK(we_N_63), 
            .Q(\mem[6] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_6__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_7__i0_i0 (.D(data[0]), .SP(we_N_63_enable_377), .CK(we_N_63), 
            .Q(\mem[7] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_7__i0_i0.GSR = "ENABLED";
    FD1P3AY mem_8__i0_i0 (.D(data[0]), .SP(we_N_63_enable_368), .CK(we_N_63), 
            .Q(\mem[8] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_8__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_9__i0_i0 (.D(data[0]), .SP(we_N_63_enable_359), .CK(we_N_63), 
            .Q(\mem[9] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_9__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_10__i0_i0 (.D(data[0]), .SP(we_N_63_enable_351), .CK(we_N_63), 
            .Q(\mem[10] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_10__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_11__i0_i0 (.D(data[0]), .SP(we_N_63_enable_343), .CK(we_N_63), 
            .Q(\mem[11] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_11__i0_i0.GSR = "ENABLED";
    FD1P3AY mem_12__i0_i0 (.D(data[0]), .SP(we_N_63_enable_336), .CK(we_N_63), 
            .Q(\mem[12] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_12__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_13__i0_i0 (.D(data[0]), .SP(we_N_63_enable_329), .CK(we_N_63), 
            .Q(\mem[13] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_13__i0_i0.GSR = "ENABLED";
    FD1P3AY mem_14__i0_i0 (.D(data[0]), .SP(we_N_63_enable_322), .CK(we_N_63), 
            .Q(\mem[14] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_14__i0_i0.GSR = "ENABLED";
    FD1P3AY mem_15__i0_i0 (.D(data[0]), .SP(we_N_63_enable_315), .CK(we_N_63), 
            .Q(\mem[15] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_15__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_16__i0_i0 (.D(data[0]), .SP(we_N_63_enable_308), .CK(we_N_63), 
            .Q(\mem[16] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_16__i0_i0.GSR = "ENABLED";
    FD1P3AY mem_17__i0_i0 (.D(data[0]), .SP(we_N_63_enable_301), .CK(we_N_63), 
            .Q(\mem[17] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_17__i0_i0.GSR = "ENABLED";
    FD1P3AY mem_18__i0_i0 (.D(data[0]), .SP(we_N_63_enable_294), .CK(we_N_63), 
            .Q(\mem[18] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_18__i0_i0.GSR = "ENABLED";
    FD1P3AY mem_19__i0_i0 (.D(data[0]), .SP(we_N_63_enable_287), .CK(we_N_63), 
            .Q(\mem[19] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_19__i0_i0.GSR = "ENABLED";
    FD1P3AY mem_20__i0_i0 (.D(data[0]), .SP(we_N_63_enable_280), .CK(we_N_63), 
            .Q(\mem[20] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_20__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_21__i0_i0 (.D(data[0]), .SP(we_N_63_enable_273), .CK(we_N_63), 
            .Q(\mem[21] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_21__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_22__i0_i0 (.D(data[0]), .SP(we_N_63_enable_266), .CK(we_N_63), 
            .Q(\mem[22] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_22__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_23__i0_i0 (.D(data[0]), .SP(we_N_63_enable_259), .CK(we_N_63), 
            .Q(\mem[23] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_23__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_24__i0_i0 (.D(data[0]), .SP(we_N_63_enable_252), .CK(we_N_63), 
            .Q(\mem[24] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_24__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_25__i0_i0 (.D(data[0]), .SP(we_N_63_enable_245), .CK(we_N_63), 
            .Q(\mem[25] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_25__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_26__i0_i0 (.D(data[0]), .SP(we_N_63_enable_238), .CK(we_N_63), 
            .Q(\mem[26] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_26__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_27__i0_i0 (.D(data[0]), .SP(we_N_63_enable_231), .CK(we_N_63), 
            .Q(\mem[27] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_27__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_28__i0_i0 (.D(data[0]), .SP(we_N_63_enable_224), .CK(we_N_63), 
            .Q(\mem[28] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_28__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_29__i0_i0 (.D(data[0]), .SP(we_N_63_enable_216), .CK(we_N_63), 
            .Q(\mem[29] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_29__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_30__i0_i0 (.D(data[0]), .SP(we_N_63_enable_201), .CK(we_N_63), 
            .Q(\mem[30] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_30__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_31__i0_i0 (.D(data[0]), .SP(we_N_63_enable_187), .CK(we_N_63), 
            .Q(\mem[31] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_31__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_32__i0_i0 (.D(data[0]), .SP(we_N_63_enable_173), .CK(we_N_63), 
            .Q(\mem[32] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_32__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_33__i0_i0 (.D(data[0]), .SP(we_N_63_enable_160), .CK(we_N_63), 
            .Q(\mem[33] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_33__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_34__i0_i0 (.D(data[0]), .SP(we_N_63_enable_129), .CK(we_N_63), 
            .Q(\mem[34] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_34__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_35__i0_i0 (.D(data[0]), .SP(we_N_63_enable_130), .CK(we_N_63), 
            .Q(\mem[35] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_35__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_36__i0_i0 (.D(data[0]), .SP(we_N_63_enable_131), .CK(we_N_63), 
            .Q(\mem[36] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_36__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_37__i0_i0 (.D(data[0]), .SP(we_N_63_enable_132), .CK(we_N_63), 
            .Q(\mem[37] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_37__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_38__i0_i0 (.D(data[0]), .SP(we_N_63_enable_133), .CK(we_N_63), 
            .Q(\mem[38] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_38__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_39__i0_i0 (.D(data[0]), .SP(we_N_63_enable_134), .CK(we_N_63), 
            .Q(\mem[39] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_39__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_40__i0_i0 (.D(data[0]), .SP(we_N_63_enable_135), .CK(we_N_63), 
            .Q(\mem[40] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_40__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_41__i0_i0 (.D(data[0]), .SP(we_N_63_enable_136), .CK(we_N_63), 
            .Q(\mem[41] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_41__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_42__i0_i0 (.D(data[0]), .SP(we_N_63_enable_137), .CK(we_N_63), 
            .Q(\mem[42] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_42__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_43__i0_i0 (.D(data[0]), .SP(we_N_63_enable_219), .CK(we_N_63), 
            .Q(\mem[43] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_43__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_44__i0_i0 (.D(data[0]), .SP(we_N_63_enable_213), .CK(we_N_63), 
            .Q(\mem[44] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_44__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_45__i0_i0 (.D(data[0]), .SP(we_N_63_enable_202), .CK(we_N_63), 
            .Q(\mem[45] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_45__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_46__i0_i0 (.D(data[0]), .SP(we_N_63_enable_188), .CK(we_N_63), 
            .Q(\mem[46] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_46__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_47__i0_i0 (.D(data[0]), .SP(we_N_63_enable_174), .CK(we_N_63), 
            .Q(\mem[47] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_47__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_48__i0_i0 (.D(data[0]), .SP(we_N_63_enable_143), .CK(we_N_63), 
            .Q(\mem[48] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_48__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_49__i0_i0 (.D(data[0]), .SP(we_N_63_enable_144), .CK(we_N_63), 
            .Q(\mem[49] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_49__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_50__i0_i0 (.D(data[0]), .SP(we_N_63_enable_512), .CK(we_N_63), 
            .Q(\mem[50] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_50__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_51__i0_i0 (.D(data[0]), .SP(we_N_63_enable_511), .CK(we_N_63), 
            .Q(\mem[51] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_51__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_52__i0_i0 (.D(data[0]), .SP(we_N_63_enable_504), .CK(we_N_63), 
            .Q(\mem[52] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_52__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_53__i0_i0 (.D(data[0]), .SP(we_N_63_enable_497), .CK(we_N_63), 
            .Q(\mem[53] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_53__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_54__i0_i0 (.D(data[0]), .SP(we_N_63_enable_490), .CK(we_N_63), 
            .Q(\mem[54] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_54__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_55__i0_i0 (.D(data[0]), .SP(we_N_63_enable_483), .CK(we_N_63), 
            .Q(\mem[55] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_55__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_56__i0_i0 (.D(data[0]), .SP(we_N_63_enable_474), .CK(we_N_63), 
            .Q(\mem[56] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_56__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_57__i0_i0 (.D(data[0]), .SP(we_N_63_enable_465), .CK(we_N_63), 
            .Q(\mem[57] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_57__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_58__i0_i0 (.D(data[0]), .SP(we_N_63_enable_455), .CK(we_N_63), 
            .Q(\mem[58] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_58__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_59__i0_i0 (.D(data[0]), .SP(we_N_63_enable_446), .CK(we_N_63), 
            .Q(\mem[59] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_59__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_60__i0_i0 (.D(data[0]), .SP(we_N_63_enable_437), .CK(we_N_63), 
            .Q(\mem[60] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_60__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_61__i0_i0 (.D(data[0]), .SP(we_N_63_enable_428), .CK(we_N_63), 
            .Q(\mem[61] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_61__i0_i0.GSR = "ENABLED";
    FD1P3AY mem_62__i0_i0 (.D(data[0]), .SP(we_N_63_enable_420), .CK(we_N_63), 
            .Q(\mem[62] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_62__i0_i0.GSR = "ENABLED";
    FD1P3AY mem_63__i0_i0 (.D(data[0]), .SP(we_N_63_enable_405), .CK(we_N_63), 
            .Q(\mem[63] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_63__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_0__i0_i0 (.D(data[0]), .SP(we_N_63_enable_379), .CK(we_N_63), 
            .Q(\mem[0] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_0__i0_i0.GSR = "ENABLED";
    FD1P3AX mem_33__i0_i1 (.D(data[1]), .SP(we_N_63_enable_160), .CK(we_N_63), 
            .Q(\mem[33] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_33__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_32__i0_i7 (.D(data[7]), .SP(we_N_63_enable_173), .CK(we_N_63), 
            .Q(\mem[32] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_32__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_47__i0_i7 (.D(data[7]), .SP(we_N_63_enable_174), .CK(we_N_63), 
            .Q(\mem[47] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_47__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_32__i0_i6 (.D(data[6]), .SP(we_N_63_enable_173), .CK(we_N_63), 
            .Q(\mem[32] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_32__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_47__i0_i6 (.D(data[6]), .SP(we_N_63_enable_174), .CK(we_N_63), 
            .Q(\mem[47] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_47__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_32__i0_i5 (.D(data[5]), .SP(we_N_63_enable_173), .CK(we_N_63), 
            .Q(\mem[32] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_32__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_47__i0_i5 (.D(data[5]), .SP(we_N_63_enable_174), .CK(we_N_63), 
            .Q(\mem[47] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_47__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_32__i0_i4 (.D(data[4]), .SP(we_N_63_enable_173), .CK(we_N_63), 
            .Q(\mem[32] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_32__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_47__i0_i4 (.D(data[4]), .SP(we_N_63_enable_174), .CK(we_N_63), 
            .Q(\mem[47] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_47__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_32__i0_i3 (.D(data[3]), .SP(we_N_63_enable_173), .CK(we_N_63), 
            .Q(\mem[32] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_32__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_47__i0_i3 (.D(data[3]), .SP(we_N_63_enable_174), .CK(we_N_63), 
            .Q(\mem[47] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_47__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_32__i0_i2 (.D(data[2]), .SP(we_N_63_enable_173), .CK(we_N_63), 
            .Q(\mem[32] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_32__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_47__i0_i2 (.D(data[2]), .SP(we_N_63_enable_174), .CK(we_N_63), 
            .Q(\mem[47] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_47__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_32__i0_i1 (.D(data[1]), .SP(we_N_63_enable_173), .CK(we_N_63), 
            .Q(\mem[32] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_32__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_47__i0_i1 (.D(data[1]), .SP(we_N_63_enable_174), .CK(we_N_63), 
            .Q(\mem[47] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_47__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_31__i0_i7 (.D(data[7]), .SP(we_N_63_enable_187), .CK(we_N_63), 
            .Q(\mem[31] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_31__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_46__i0_i7 (.D(data[7]), .SP(we_N_63_enable_188), .CK(we_N_63), 
            .Q(\mem[46] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_46__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_31__i0_i6 (.D(data[6]), .SP(we_N_63_enable_187), .CK(we_N_63), 
            .Q(\mem[31] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_31__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_46__i0_i6 (.D(data[6]), .SP(we_N_63_enable_188), .CK(we_N_63), 
            .Q(\mem[46] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_46__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_31__i0_i5 (.D(data[5]), .SP(we_N_63_enable_187), .CK(we_N_63), 
            .Q(\mem[31] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_31__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_46__i0_i5 (.D(data[5]), .SP(we_N_63_enable_188), .CK(we_N_63), 
            .Q(\mem[46] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_46__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_31__i0_i4 (.D(data[4]), .SP(we_N_63_enable_187), .CK(we_N_63), 
            .Q(\mem[31] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_31__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_46__i0_i4 (.D(data[4]), .SP(we_N_63_enable_188), .CK(we_N_63), 
            .Q(\mem[46] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_46__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_31__i0_i3 (.D(data[3]), .SP(we_N_63_enable_187), .CK(we_N_63), 
            .Q(\mem[31] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_31__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_46__i0_i3 (.D(data[3]), .SP(we_N_63_enable_188), .CK(we_N_63), 
            .Q(\mem[46] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_46__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_31__i0_i2 (.D(data[2]), .SP(we_N_63_enable_187), .CK(we_N_63), 
            .Q(\mem[31] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_31__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_46__i0_i2 (.D(data[2]), .SP(we_N_63_enable_188), .CK(we_N_63), 
            .Q(\mem[46] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_46__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_31__i0_i1 (.D(data[1]), .SP(we_N_63_enable_187), .CK(we_N_63), 
            .Q(\mem[31] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_31__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_46__i0_i1 (.D(data[1]), .SP(we_N_63_enable_188), .CK(we_N_63), 
            .Q(\mem[46] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_46__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_30__i0_i7 (.D(data[7]), .SP(we_N_63_enable_201), .CK(we_N_63), 
            .Q(\mem[30] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_30__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_45__i0_i7 (.D(data[7]), .SP(we_N_63_enable_202), .CK(we_N_63), 
            .Q(\mem[45] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_45__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_30__i0_i6 (.D(data[6]), .SP(we_N_63_enable_201), .CK(we_N_63), 
            .Q(\mem[30] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_30__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_45__i0_i6 (.D(data[6]), .SP(we_N_63_enable_202), .CK(we_N_63), 
            .Q(\mem[45] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_45__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_30__i0_i5 (.D(data[5]), .SP(we_N_63_enable_201), .CK(we_N_63), 
            .Q(\mem[30] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_30__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_45__i0_i5 (.D(data[5]), .SP(we_N_63_enable_202), .CK(we_N_63), 
            .Q(\mem[45] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_45__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_30__i0_i4 (.D(data[4]), .SP(we_N_63_enable_201), .CK(we_N_63), 
            .Q(\mem[30] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_30__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_45__i0_i4 (.D(data[4]), .SP(we_N_63_enable_202), .CK(we_N_63), 
            .Q(\mem[45] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_45__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_30__i0_i3 (.D(data[3]), .SP(we_N_63_enable_201), .CK(we_N_63), 
            .Q(\mem[30] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_30__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_45__i0_i3 (.D(data[3]), .SP(we_N_63_enable_202), .CK(we_N_63), 
            .Q(\mem[45] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_45__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_30__i0_i2 (.D(data[2]), .SP(we_N_63_enable_201), .CK(we_N_63), 
            .Q(\mem[30] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_30__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_45__i0_i2 (.D(data[2]), .SP(we_N_63_enable_202), .CK(we_N_63), 
            .Q(\mem[45] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_45__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_30__i0_i1 (.D(data[1]), .SP(we_N_63_enable_201), .CK(we_N_63), 
            .Q(\mem[30] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_30__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_45__i0_i1 (.D(data[1]), .SP(we_N_63_enable_202), .CK(we_N_63), 
            .Q(\mem[45] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_45__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_29__i0_i7 (.D(data[7]), .SP(we_N_63_enable_216), .CK(we_N_63), 
            .Q(\mem[29] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_29__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_44__i0_i7 (.D(data[7]), .SP(we_N_63_enable_213), .CK(we_N_63), 
            .Q(\mem[44] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_44__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_29__i0_i6 (.D(data[6]), .SP(we_N_63_enable_216), .CK(we_N_63), 
            .Q(\mem[29] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_29__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_44__i0_i6 (.D(data[6]), .SP(we_N_63_enable_213), .CK(we_N_63), 
            .Q(\mem[44] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_44__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_29__i0_i5 (.D(data[5]), .SP(we_N_63_enable_216), .CK(we_N_63), 
            .Q(\mem[29] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_29__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_44__i0_i5 (.D(data[5]), .SP(we_N_63_enable_213), .CK(we_N_63), 
            .Q(\mem[44] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_44__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_29__i0_i4 (.D(data[4]), .SP(we_N_63_enable_216), .CK(we_N_63), 
            .Q(\mem[29] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_29__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_44__i0_i4 (.D(data[4]), .SP(we_N_63_enable_213), .CK(we_N_63), 
            .Q(\mem[44] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_44__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_44__i0_i3 (.D(data[3]), .SP(we_N_63_enable_213), .CK(we_N_63), 
            .Q(\mem[44] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_44__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_44__i0_i2 (.D(data[2]), .SP(we_N_63_enable_213), .CK(we_N_63), 
            .Q(\mem[44] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_44__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_44__i0_i1 (.D(data[1]), .SP(we_N_63_enable_213), .CK(we_N_63), 
            .Q(\mem[44] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_44__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_29__i0_i3 (.D(data[3]), .SP(we_N_63_enable_216), .CK(we_N_63), 
            .Q(\mem[29] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_29__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_29__i0_i2 (.D(data[2]), .SP(we_N_63_enable_216), .CK(we_N_63), 
            .Q(\mem[29] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_29__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_29__i0_i1 (.D(data[1]), .SP(we_N_63_enable_216), .CK(we_N_63), 
            .Q(\mem[29] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_29__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_28__i0_i7 (.D(data[7]), .SP(we_N_63_enable_224), .CK(we_N_63), 
            .Q(\mem[28] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_28__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_28__i0_i6 (.D(data[6]), .SP(we_N_63_enable_224), .CK(we_N_63), 
            .Q(\mem[28] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_28__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_43__i0_i7 (.D(data[7]), .SP(we_N_63_enable_219), .CK(we_N_63), 
            .Q(\mem[43] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_43__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_28__i0_i5 (.D(data[5]), .SP(we_N_63_enable_224), .CK(we_N_63), 
            .Q(\mem[28] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_28__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_28__i0_i4 (.D(data[4]), .SP(we_N_63_enable_224), .CK(we_N_63), 
            .Q(\mem[28] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_28__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_28__i0_i3 (.D(data[3]), .SP(we_N_63_enable_224), .CK(we_N_63), 
            .Q(\mem[28] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_28__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_28__i0_i2 (.D(data[2]), .SP(we_N_63_enable_224), .CK(we_N_63), 
            .Q(\mem[28] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_28__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_28__i0_i1 (.D(data[1]), .SP(we_N_63_enable_224), .CK(we_N_63), 
            .Q(\mem[28] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_28__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_27__i0_i7 (.D(data[7]), .SP(we_N_63_enable_231), .CK(we_N_63), 
            .Q(\mem[27] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_27__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_27__i0_i6 (.D(data[6]), .SP(we_N_63_enable_231), .CK(we_N_63), 
            .Q(\mem[27] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_27__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_27__i0_i5 (.D(data[5]), .SP(we_N_63_enable_231), .CK(we_N_63), 
            .Q(\mem[27] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_27__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_27__i0_i4 (.D(data[4]), .SP(we_N_63_enable_231), .CK(we_N_63), 
            .Q(\mem[27] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_27__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_27__i0_i3 (.D(data[3]), .SP(we_N_63_enable_231), .CK(we_N_63), 
            .Q(\mem[27] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_27__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_27__i0_i2 (.D(data[2]), .SP(we_N_63_enable_231), .CK(we_N_63), 
            .Q(\mem[27] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_27__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_27__i0_i1 (.D(data[1]), .SP(we_N_63_enable_231), .CK(we_N_63), 
            .Q(\mem[27] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_27__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_26__i0_i7 (.D(data[7]), .SP(we_N_63_enable_238), .CK(we_N_63), 
            .Q(\mem[26] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_26__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_26__i0_i6 (.D(data[6]), .SP(we_N_63_enable_238), .CK(we_N_63), 
            .Q(\mem[26] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_26__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_26__i0_i5 (.D(data[5]), .SP(we_N_63_enable_238), .CK(we_N_63), 
            .Q(\mem[26] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_26__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_26__i0_i4 (.D(data[4]), .SP(we_N_63_enable_238), .CK(we_N_63), 
            .Q(\mem[26] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_26__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_26__i0_i3 (.D(data[3]), .SP(we_N_63_enable_238), .CK(we_N_63), 
            .Q(\mem[26] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_26__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_26__i0_i2 (.D(data[2]), .SP(we_N_63_enable_238), .CK(we_N_63), 
            .Q(\mem[26] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_26__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_26__i0_i1 (.D(data[1]), .SP(we_N_63_enable_238), .CK(we_N_63), 
            .Q(\mem[26] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_26__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_25__i0_i7 (.D(data[7]), .SP(we_N_63_enable_245), .CK(we_N_63), 
            .Q(\mem[25] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_25__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_25__i0_i6 (.D(data[6]), .SP(we_N_63_enable_245), .CK(we_N_63), 
            .Q(\mem[25] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_25__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_25__i0_i5 (.D(data[5]), .SP(we_N_63_enable_245), .CK(we_N_63), 
            .Q(\mem[25] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_25__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_25__i0_i4 (.D(data[4]), .SP(we_N_63_enable_245), .CK(we_N_63), 
            .Q(\mem[25] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_25__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_25__i0_i3 (.D(data[3]), .SP(we_N_63_enable_245), .CK(we_N_63), 
            .Q(\mem[25] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_25__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_25__i0_i2 (.D(data[2]), .SP(we_N_63_enable_245), .CK(we_N_63), 
            .Q(\mem[25] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_25__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_25__i0_i1 (.D(data[1]), .SP(we_N_63_enable_245), .CK(we_N_63), 
            .Q(\mem[25] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_25__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_24__i0_i7 (.D(data[7]), .SP(we_N_63_enable_252), .CK(we_N_63), 
            .Q(\mem[24] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_24__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_24__i0_i6 (.D(data[6]), .SP(we_N_63_enable_252), .CK(we_N_63), 
            .Q(\mem[24] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_24__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_24__i0_i5 (.D(data[5]), .SP(we_N_63_enable_252), .CK(we_N_63), 
            .Q(\mem[24] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_24__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_24__i0_i4 (.D(data[4]), .SP(we_N_63_enable_252), .CK(we_N_63), 
            .Q(\mem[24] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_24__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_24__i0_i3 (.D(data[3]), .SP(we_N_63_enable_252), .CK(we_N_63), 
            .Q(\mem[24] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_24__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_24__i0_i2 (.D(data[2]), .SP(we_N_63_enable_252), .CK(we_N_63), 
            .Q(\mem[24] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_24__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_24__i0_i1 (.D(data[1]), .SP(we_N_63_enable_252), .CK(we_N_63), 
            .Q(\mem[24] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_24__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_23__i0_i7 (.D(data[7]), .SP(we_N_63_enable_259), .CK(we_N_63), 
            .Q(\mem[23] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_23__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_23__i0_i6 (.D(data[6]), .SP(we_N_63_enable_259), .CK(we_N_63), 
            .Q(\mem[23] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_23__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_23__i0_i5 (.D(data[5]), .SP(we_N_63_enable_259), .CK(we_N_63), 
            .Q(\mem[23] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_23__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_23__i0_i4 (.D(data[4]), .SP(we_N_63_enable_259), .CK(we_N_63), 
            .Q(\mem[23] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_23__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_23__i0_i3 (.D(data[3]), .SP(we_N_63_enable_259), .CK(we_N_63), 
            .Q(\mem[23] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_23__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_23__i0_i2 (.D(data[2]), .SP(we_N_63_enable_259), .CK(we_N_63), 
            .Q(\mem[23] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_23__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_23__i0_i1 (.D(data[1]), .SP(we_N_63_enable_259), .CK(we_N_63), 
            .Q(\mem[23] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_23__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_22__i0_i7 (.D(data[7]), .SP(we_N_63_enable_266), .CK(we_N_63), 
            .Q(\mem[22] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_22__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_22__i0_i6 (.D(data[6]), .SP(we_N_63_enable_266), .CK(we_N_63), 
            .Q(\mem[22] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_22__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_22__i0_i5 (.D(data[5]), .SP(we_N_63_enable_266), .CK(we_N_63), 
            .Q(\mem[22] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_22__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_22__i0_i4 (.D(data[4]), .SP(we_N_63_enable_266), .CK(we_N_63), 
            .Q(\mem[22] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_22__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_22__i0_i3 (.D(data[3]), .SP(we_N_63_enable_266), .CK(we_N_63), 
            .Q(\mem[22] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_22__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_22__i0_i2 (.D(data[2]), .SP(we_N_63_enable_266), .CK(we_N_63), 
            .Q(\mem[22] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_22__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_22__i0_i1 (.D(data[1]), .SP(we_N_63_enable_266), .CK(we_N_63), 
            .Q(\mem[22] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_22__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_21__i0_i7 (.D(data[7]), .SP(we_N_63_enable_273), .CK(we_N_63), 
            .Q(\mem[21] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_21__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_21__i0_i6 (.D(data[6]), .SP(we_N_63_enable_273), .CK(we_N_63), 
            .Q(\mem[21] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_21__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_21__i0_i5 (.D(data[5]), .SP(we_N_63_enable_273), .CK(we_N_63), 
            .Q(\mem[21] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_21__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_21__i0_i4 (.D(data[4]), .SP(we_N_63_enable_273), .CK(we_N_63), 
            .Q(\mem[21] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_21__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_21__i0_i3 (.D(data[3]), .SP(we_N_63_enable_273), .CK(we_N_63), 
            .Q(\mem[21] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_21__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_21__i0_i2 (.D(data[2]), .SP(we_N_63_enable_273), .CK(we_N_63), 
            .Q(\mem[21] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_21__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_21__i0_i1 (.D(data[1]), .SP(we_N_63_enable_273), .CK(we_N_63), 
            .Q(\mem[21] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_21__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_20__i0_i7 (.D(data[7]), .SP(we_N_63_enable_280), .CK(we_N_63), 
            .Q(\mem[20] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_20__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_20__i0_i6 (.D(data[6]), .SP(we_N_63_enable_280), .CK(we_N_63), 
            .Q(\mem[20] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_20__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_20__i0_i5 (.D(data[5]), .SP(we_N_63_enable_280), .CK(we_N_63), 
            .Q(\mem[20] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_20__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_20__i0_i4 (.D(data[4]), .SP(we_N_63_enable_280), .CK(we_N_63), 
            .Q(\mem[20] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_20__i0_i4.GSR = "ENABLED";
    FD1P3AY mem_20__i0_i3 (.D(data[3]), .SP(we_N_63_enable_280), .CK(we_N_63), 
            .Q(\mem[20] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_20__i0_i3.GSR = "ENABLED";
    FD1P3AY mem_20__i0_i2 (.D(data[2]), .SP(we_N_63_enable_280), .CK(we_N_63), 
            .Q(\mem[20] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_20__i0_i2.GSR = "ENABLED";
    FD1P3AY mem_20__i0_i1 (.D(data[1]), .SP(we_N_63_enable_280), .CK(we_N_63), 
            .Q(\mem[20] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_20__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_19__i0_i7 (.D(data[7]), .SP(we_N_63_enable_287), .CK(we_N_63), 
            .Q(\mem[19] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_19__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_19__i0_i6 (.D(data[6]), .SP(we_N_63_enable_287), .CK(we_N_63), 
            .Q(\mem[19] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_19__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_19__i0_i5 (.D(data[5]), .SP(we_N_63_enable_287), .CK(we_N_63), 
            .Q(\mem[19] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_19__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_19__i0_i4 (.D(data[4]), .SP(we_N_63_enable_287), .CK(we_N_63), 
            .Q(\mem[19] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_19__i0_i4.GSR = "ENABLED";
    FD1P3AY mem_19__i0_i3 (.D(data[3]), .SP(we_N_63_enable_287), .CK(we_N_63), 
            .Q(\mem[19] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_19__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_19__i0_i2 (.D(data[2]), .SP(we_N_63_enable_287), .CK(we_N_63), 
            .Q(\mem[19] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_19__i0_i2.GSR = "ENABLED";
    LUT4 Select_676_i3_4_lut (.A(data_7__N_66[0]), .B(akku_o_c_0), .C(oe_N_57), 
         .D(n2305), .Z(data[0])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((D)+!B)) */ ;
    defparam Select_676_i3_4_lut.init = 16'ha0ec;
    FD1P3AX mem_19__i0_i1 (.D(data[1]), .SP(we_N_63_enable_287), .CK(we_N_63), 
            .Q(\mem[19] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_19__i0_i1.GSR = "ENABLED";
    LUT4 Select_671_i3_4_lut (.A(data_7__N_66[5]), .B(akku_o_c_5), .C(oe_N_57), 
         .D(n2305), .Z(data[5])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((D)+!B)) */ ;
    defparam Select_671_i3_4_lut.init = 16'ha0ec;
    FD1P3AY mem_18__i0_i7 (.D(data[7]), .SP(we_N_63_enable_294), .CK(we_N_63), 
            .Q(\mem[18] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_18__i0_i7.GSR = "ENABLED";
    FD1P3AY mem_18__i0_i6 (.D(data[6]), .SP(we_N_63_enable_294), .CK(we_N_63), 
            .Q(\mem[18] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_18__i0_i6.GSR = "ENABLED";
    LUT4 i1771_3_lut (.A(\mem[38] [5]), .B(\mem[39] [5]), .C(\adrram[0] ), 
         .Z(n1904)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1771_3_lut.init = 16'hcaca;
    FD1P3AX mem_18__i0_i5 (.D(data[5]), .SP(we_N_63_enable_294), .CK(we_N_63), 
            .Q(\mem[18] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_18__i0_i5.GSR = "ENABLED";
    FD1P3AY mem_18__i0_i4 (.D(data[4]), .SP(we_N_63_enable_294), .CK(we_N_63), 
            .Q(\mem[18] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_18__i0_i4.GSR = "ENABLED";
    LUT4 i1770_3_lut (.A(\mem[36] [5]), .B(\mem[37] [5]), .C(\adrram[0] ), 
         .Z(n1903)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1770_3_lut.init = 16'hcaca;
    LUT4 i1872_3_lut (.A(\mem[54] [2]), .B(\mem[55] [2]), .C(\adrram[0] ), 
         .Z(n2005)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1872_3_lut.init = 16'hcaca;
    FD1P3AX mem_18__i0_i3 (.D(data[3]), .SP(we_N_63_enable_294), .CK(we_N_63), 
            .Q(\mem[18] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_18__i0_i3.GSR = "ENABLED";
    LUT4 i1871_3_lut (.A(\mem[52] [2]), .B(\mem[53] [2]), .C(\adrram[0] ), 
         .Z(n2004)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1871_3_lut.init = 16'hcaca;
    FD1P3AX mem_18__i0_i2 (.D(data[2]), .SP(we_N_63_enable_294), .CK(we_N_63), 
            .Q(\mem[18] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_18__i0_i2.GSR = "ENABLED";
    LUT4 i1769_3_lut (.A(\mem[34] [5]), .B(\mem[35] [5]), .C(\adrram[0] ), 
         .Z(n1902)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1769_3_lut.init = 16'hcaca;
    FD1P3AX mem_18__i0_i1 (.D(data[1]), .SP(we_N_63_enable_294), .CK(we_N_63), 
            .Q(\mem[18] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_18__i0_i1.GSR = "ENABLED";
    FD1P3AY mem_17__i0_i7 (.D(data[7]), .SP(we_N_63_enable_301), .CK(we_N_63), 
            .Q(\mem[17] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_17__i0_i7.GSR = "ENABLED";
    FD1P3AY mem_17__i0_i6 (.D(data[6]), .SP(we_N_63_enable_301), .CK(we_N_63), 
            .Q(\mem[17] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_17__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_17__i0_i5 (.D(data[5]), .SP(we_N_63_enable_301), .CK(we_N_63), 
            .Q(\mem[17] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_17__i0_i5.GSR = "ENABLED";
    LUT4 i1768_3_lut (.A(\mem[32] [5]), .B(\mem[33] [5]), .C(\adrram[0] ), 
         .Z(n1901)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1768_3_lut.init = 16'hcaca;
    LUT4 i1870_3_lut (.A(\mem[50] [2]), .B(\mem[51] [2]), .C(\adrram[0] ), 
         .Z(n2003)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1870_3_lut.init = 16'hcaca;
    FD1P3AY mem_17__i0_i4 (.D(data[4]), .SP(we_N_63_enable_301), .CK(we_N_63), 
            .Q(\mem[17] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_17__i0_i4.GSR = "ENABLED";
    LUT4 i1869_3_lut (.A(\mem[48] [2]), .B(\mem[49] [2]), .C(\adrram[0] ), 
         .Z(n2002)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1869_3_lut.init = 16'hcaca;
    FD1P3AX mem_17__i0_i3 (.D(data[3]), .SP(we_N_63_enable_301), .CK(we_N_63), 
            .Q(\mem[17] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_17__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_17__i0_i2 (.D(data[2]), .SP(we_N_63_enable_301), .CK(we_N_63), 
            .Q(\mem[17] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_17__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_17__i0_i1 (.D(data[1]), .SP(we_N_63_enable_301), .CK(we_N_63), 
            .Q(\mem[17] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_17__i0_i1.GSR = "ENABLED";
    FD1P3AY mem_16__i0_i7 (.D(data[7]), .SP(we_N_63_enable_308), .CK(we_N_63), 
            .Q(\mem[16] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_16__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_16__i0_i6 (.D(data[6]), .SP(we_N_63_enable_308), .CK(we_N_63), 
            .Q(\mem[16] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_16__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_16__i0_i5 (.D(data[5]), .SP(we_N_63_enable_308), .CK(we_N_63), 
            .Q(\mem[16] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_16__i0_i5.GSR = "ENABLED";
    LUT4 i1868_3_lut (.A(\mem[46] [2]), .B(\mem[47] [2]), .C(\adrram[0] ), 
         .Z(n2001)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1868_3_lut.init = 16'hcaca;
    FD1P3AY mem_16__i0_i4 (.D(data[4]), .SP(we_N_63_enable_308), .CK(we_N_63), 
            .Q(\mem[16] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_16__i0_i4.GSR = "ENABLED";
    LUT4 i1867_3_lut (.A(\mem[44] [2]), .B(\mem[45] [2]), .C(\adrram[0] ), 
         .Z(n2000)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1867_3_lut.init = 16'hcaca;
    FD1P3AX mem_16__i0_i3 (.D(data[3]), .SP(we_N_63_enable_308), .CK(we_N_63), 
            .Q(\mem[16] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_16__i0_i3.GSR = "ENABLED";
    FD1P3AY mem_16__i0_i2 (.D(data[2]), .SP(we_N_63_enable_308), .CK(we_N_63), 
            .Q(\mem[16] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_16__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_16__i0_i1 (.D(data[1]), .SP(we_N_63_enable_308), .CK(we_N_63), 
            .Q(\mem[16] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_16__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_15__i0_i7 (.D(data[7]), .SP(we_N_63_enable_315), .CK(we_N_63), 
            .Q(\mem[15] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_15__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_15__i0_i6 (.D(data[6]), .SP(we_N_63_enable_315), .CK(we_N_63), 
            .Q(\mem[15] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_15__i0_i6.GSR = "ENABLED";
    LUT4 i1866_3_lut (.A(\mem[42] [2]), .B(\mem[43] [2]), .C(\adrram[0] ), 
         .Z(n1999)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1866_3_lut.init = 16'hcaca;
    FD1P3AY mem_15__i0_i5 (.D(data[5]), .SP(we_N_63_enable_315), .CK(we_N_63), 
            .Q(\mem[15] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_15__i0_i5.GSR = "ENABLED";
    LUT4 i1865_3_lut (.A(\mem[40] [2]), .B(\mem[41] [2]), .C(\adrram[0] ), 
         .Z(n1998)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1865_3_lut.init = 16'hcaca;
    FD1P3AY mem_15__i0_i4 (.D(data[4]), .SP(we_N_63_enable_315), .CK(we_N_63), 
            .Q(\mem[15] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_15__i0_i4.GSR = "ENABLED";
    LUT4 i1469_3_lut (.A(\mem[22] [0]), .B(\mem[23] [0]), .C(\adrram[0] ), 
         .Z(n1602)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1469_3_lut.init = 16'hcaca;
    FD1P3AY mem_15__i0_i3 (.D(data[3]), .SP(we_N_63_enable_315), .CK(we_N_63), 
            .Q(\mem[15] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_15__i0_i3.GSR = "ENABLED";
    FD1P3AY mem_15__i0_i2 (.D(data[2]), .SP(we_N_63_enable_315), .CK(we_N_63), 
            .Q(\mem[15] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_15__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_15__i0_i1 (.D(data[1]), .SP(we_N_63_enable_315), .CK(we_N_63), 
            .Q(\mem[15] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_15__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_14__i0_i7 (.D(data[7]), .SP(we_N_63_enable_322), .CK(we_N_63), 
            .Q(\mem[14] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_14__i0_i7.GSR = "ENABLED";
    LUT4 i1468_3_lut (.A(\mem[20] [0]), .B(\mem[21] [0]), .C(\adrram[0] ), 
         .Z(n1601)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1468_3_lut.init = 16'hcaca;
    FD1P3AY mem_14__i0_i6 (.D(data[6]), .SP(we_N_63_enable_322), .CK(we_N_63), 
            .Q(\mem[14] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_14__i0_i6.GSR = "ENABLED";
    LUT4 i1864_3_lut (.A(\mem[38] [2]), .B(\mem[39] [2]), .C(\adrram[0] ), 
         .Z(n1997)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1864_3_lut.init = 16'hcaca;
    FD1P3AX mem_14__i0_i5 (.D(data[5]), .SP(we_N_63_enable_322), .CK(we_N_63), 
            .Q(\mem[14] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_14__i0_i5.GSR = "ENABLED";
    LUT4 i1863_3_lut (.A(\mem[36] [2]), .B(\mem[37] [2]), .C(\adrram[0] ), 
         .Z(n1996)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1863_3_lut.init = 16'hcaca;
    FD1P3AY mem_14__i0_i4 (.D(data[4]), .SP(we_N_63_enable_322), .CK(we_N_63), 
            .Q(\mem[14] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_14__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_14__i0_i3 (.D(data[3]), .SP(we_N_63_enable_322), .CK(we_N_63), 
            .Q(\mem[14] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_14__i0_i3.GSR = "ENABLED";
    FD1P3AY mem_14__i0_i2 (.D(data[2]), .SP(we_N_63_enable_322), .CK(we_N_63), 
            .Q(\mem[14] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_14__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_14__i0_i1 (.D(data[1]), .SP(we_N_63_enable_322), .CK(we_N_63), 
            .Q(\mem[14] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_14__i0_i1.GSR = "ENABLED";
    LUT4 i1862_3_lut (.A(\mem[34] [2]), .B(\mem[35] [2]), .C(\adrram[0] ), 
         .Z(n1995)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1862_3_lut.init = 16'hcaca;
    FD1P3AY mem_13__i0_i7 (.D(data[7]), .SP(we_N_63_enable_329), .CK(we_N_63), 
            .Q(\mem[13] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_13__i0_i7.GSR = "ENABLED";
    LUT4 i1861_3_lut (.A(\mem[32] [2]), .B(\mem[33] [2]), .C(\adrram[0] ), 
         .Z(n1994)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1861_3_lut.init = 16'hcaca;
    LUT4 i1467_3_lut (.A(\mem[18] [0]), .B(\mem[19] [0]), .C(\adrram[0] ), 
         .Z(n1600)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1467_3_lut.init = 16'hcaca;
    FD1P3AY mem_13__i0_i6 (.D(data[6]), .SP(we_N_63_enable_329), .CK(we_N_63), 
            .Q(\mem[13] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_13__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_13__i0_i5 (.D(data[5]), .SP(we_N_63_enable_329), .CK(we_N_63), 
            .Q(\mem[13] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_13__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_13__i0_i4 (.D(data[4]), .SP(we_N_63_enable_329), .CK(we_N_63), 
            .Q(\mem[13] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_13__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_13__i0_i3 (.D(data[3]), .SP(we_N_63_enable_329), .CK(we_N_63), 
            .Q(\mem[13] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_13__i0_i3.GSR = "ENABLED";
    FD1P3AY mem_13__i0_i2 (.D(data[2]), .SP(we_N_63_enable_329), .CK(we_N_63), 
            .Q(\mem[13] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_13__i0_i2.GSR = "ENABLED";
    FD1P3AY mem_13__i0_i1 (.D(data[1]), .SP(we_N_63_enable_329), .CK(we_N_63), 
            .Q(\mem[13] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_13__i0_i1.GSR = "ENABLED";
    LUT4 i1466_3_lut (.A(\mem[16] [0]), .B(\mem[17] [0]), .C(\adrram[0] ), 
         .Z(n1599)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1466_3_lut.init = 16'hcaca;
    FD1P3AY mem_12__i0_i7 (.D(data[7]), .SP(we_N_63_enable_336), .CK(we_N_63), 
            .Q(\mem[12] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_12__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_12__i0_i6 (.D(data[6]), .SP(we_N_63_enable_336), .CK(we_N_63), 
            .Q(\mem[12] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_12__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_12__i0_i5 (.D(data[5]), .SP(we_N_63_enable_336), .CK(we_N_63), 
            .Q(\mem[12] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_12__i0_i5.GSR = "ENABLED";
    FD1P3AY mem_12__i0_i4 (.D(data[4]), .SP(we_N_63_enable_336), .CK(we_N_63), 
            .Q(\mem[12] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_12__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_12__i0_i3 (.D(data[3]), .SP(we_N_63_enable_336), .CK(we_N_63), 
            .Q(\mem[12] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_12__i0_i3.GSR = "ENABLED";
    FD1P3AY mem_12__i0_i2 (.D(data[2]), .SP(we_N_63_enable_336), .CK(we_N_63), 
            .Q(\mem[12] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_12__i0_i2.GSR = "ENABLED";
    LUT4 i1465_3_lut (.A(\mem[14] [0]), .B(\mem[15] [0]), .C(\adrram[0] ), 
         .Z(n1598)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1465_3_lut.init = 16'hcaca;
    FD1P3AX mem_12__i0_i1 (.D(data[1]), .SP(we_N_63_enable_336), .CK(we_N_63), 
            .Q(\mem[12] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_12__i0_i1.GSR = "ENABLED";
    FD1P3AY mem_11__i0_i7 (.D(data[7]), .SP(we_N_63_enable_343), .CK(we_N_63), 
            .Q(\mem[11] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_11__i0_i7.GSR = "ENABLED";
    FD1P3AY mem_11__i0_i6 (.D(data[6]), .SP(we_N_63_enable_343), .CK(we_N_63), 
            .Q(\mem[11] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_11__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_11__i0_i5 (.D(data[5]), .SP(we_N_63_enable_343), .CK(we_N_63), 
            .Q(\mem[11] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_11__i0_i5.GSR = "ENABLED";
    LUT4 i1464_3_lut (.A(\mem[12] [0]), .B(\mem[13] [0]), .C(\adrram[0] ), 
         .Z(n1597)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1464_3_lut.init = 16'hcaca;
    FD1P3AX mem_11__i0_i4 (.D(data[4]), .SP(we_N_63_enable_343), .CK(we_N_63), 
            .Q(\mem[11] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_11__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_11__i0_i3 (.D(data[3]), .SP(we_N_63_enable_343), .CK(we_N_63), 
            .Q(\mem[11] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_11__i0_i3.GSR = "ENABLED";
    FD1P3AY mem_11__i0_i2 (.D(data[2]), .SP(we_N_63_enable_343), .CK(we_N_63), 
            .Q(\mem[11] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_11__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_11__i0_i1 (.D(data[1]), .SP(we_N_63_enable_343), .CK(we_N_63), 
            .Q(\mem[11] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_11__i0_i1.GSR = "ENABLED";
    FD1P3AY mem_10__i0_i7 (.D(data[7]), .SP(we_N_63_enable_351), .CK(we_N_63), 
            .Q(\mem[10] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_10__i0_i7.GSR = "ENABLED";
    LUT4 i1463_3_lut (.A(\mem[10] [0]), .B(\mem[11] [0]), .C(\adrram[0] ), 
         .Z(n1596)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1463_3_lut.init = 16'hcaca;
    FD1P3AX mem_0__i0_i7 (.D(data[7]), .SP(we_N_63_enable_379), .CK(we_N_63), 
            .Q(\mem[0] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_0__i0_i7.GSR = "ENABLED";
    FD1P3AY mem_10__i0_i6 (.D(data[6]), .SP(we_N_63_enable_351), .CK(we_N_63), 
            .Q(\mem[10] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_10__i0_i6.GSR = "ENABLED";
    LUT4 i1462_3_lut (.A(\mem[8] [0]), .B(\mem[9] [0]), .C(\adrram[0] ), 
         .Z(n1595)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1462_3_lut.init = 16'hcaca;
    FD1P3AX mem_10__i0_i5 (.D(data[5]), .SP(we_N_63_enable_351), .CK(we_N_63), 
            .Q(\mem[10] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_10__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_10__i0_i4 (.D(data[4]), .SP(we_N_63_enable_351), .CK(we_N_63), 
            .Q(\mem[10] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_10__i0_i4.GSR = "ENABLED";
    FD1P3AY mem_10__i0_i3 (.D(data[3]), .SP(we_N_63_enable_351), .CK(we_N_63), 
            .Q(\mem[10] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_10__i0_i3.GSR = "ENABLED";
    FD1P3AY mem_10__i0_i2 (.D(data[2]), .SP(we_N_63_enable_351), .CK(we_N_63), 
            .Q(\mem[10] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_10__i0_i2.GSR = "ENABLED";
    FD1P3AY mem_10__i0_i1 (.D(data[1]), .SP(we_N_63_enable_351), .CK(we_N_63), 
            .Q(\mem[10] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_10__i0_i1.GSR = "ENABLED";
    LUT4 i1566_3_lut (.A(\mem[30] [3]), .B(\mem[31] [3]), .C(\adrram[0] ), 
         .Z(n1699)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1566_3_lut.init = 16'hcaca;
    FD1P3AX mem_9__i0_i7 (.D(data[7]), .SP(we_N_63_enable_359), .CK(we_N_63), 
            .Q(\mem[9] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_9__i0_i7.GSR = "ENABLED";
    FD1P3AY mem_9__i0_i6 (.D(data[6]), .SP(we_N_63_enable_359), .CK(we_N_63), 
            .Q(\mem[9] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_9__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_0__i0_i6 (.D(data[6]), .SP(we_N_63_enable_379), .CK(we_N_63), 
            .Q(\mem[0] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_0__i0_i6.GSR = "ENABLED";
    FD1P3AY mem_9__i0_i5 (.D(data[5]), .SP(we_N_63_enable_359), .CK(we_N_63), 
            .Q(\mem[9] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_9__i0_i5.GSR = "ENABLED";
    FD1P3AY mem_9__i0_i4 (.D(data[4]), .SP(we_N_63_enable_359), .CK(we_N_63), 
            .Q(\mem[9] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_9__i0_i4.GSR = "ENABLED";
    FD1P3AY mem_9__i0_i3 (.D(data[3]), .SP(we_N_63_enable_359), .CK(we_N_63), 
            .Q(\mem[9] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_9__i0_i3.GSR = "ENABLED";
    FD1P3AY mem_9__i0_i2 (.D(data[2]), .SP(we_N_63_enable_359), .CK(we_N_63), 
            .Q(\mem[9] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_9__i0_i2.GSR = "ENABLED";
    FD1P3AY mem_9__i0_i1 (.D(data[1]), .SP(we_N_63_enable_359), .CK(we_N_63), 
            .Q(\mem[9] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_9__i0_i1.GSR = "ENABLED";
    FD1P3AY mem_8__i0_i7 (.D(data[7]), .SP(we_N_63_enable_368), .CK(we_N_63), 
            .Q(\mem[8] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_8__i0_i7.GSR = "ENABLED";
    LUT4 i1565_3_lut (.A(\mem[28] [3]), .B(\mem[29] [3]), .C(\adrram[0] ), 
         .Z(n1698)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1565_3_lut.init = 16'hcaca;
    FD1P3AX mem_8__i0_i6 (.D(data[6]), .SP(we_N_63_enable_368), .CK(we_N_63), 
            .Q(\mem[8] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_8__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_8__i0_i5 (.D(data[5]), .SP(we_N_63_enable_368), .CK(we_N_63), 
            .Q(\mem[8] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_8__i0_i5.GSR = "ENABLED";
    FD1P3AY mem_0__i0_i5 (.D(data[5]), .SP(we_N_63_enable_379), .CK(we_N_63), 
            .Q(\mem[0] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_0__i0_i5.GSR = "ENABLED";
    FD1P3AY mem_0__i0_i4 (.D(data[4]), .SP(we_N_63_enable_379), .CK(we_N_63), 
            .Q(\mem[0] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_0__i0_i4.GSR = "ENABLED";
    FD1P3AY mem_8__i0_i4 (.D(data[4]), .SP(we_N_63_enable_368), .CK(we_N_63), 
            .Q(\mem[8] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_8__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_8__i0_i3 (.D(data[3]), .SP(we_N_63_enable_368), .CK(we_N_63), 
            .Q(\mem[8] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_8__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_8__i0_i2 (.D(data[2]), .SP(we_N_63_enable_368), .CK(we_N_63), 
            .Q(\mem[8] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_8__i0_i2.GSR = "ENABLED";
    LUT4 i1461_3_lut (.A(\mem[6] [0]), .B(\mem[7] [0]), .C(\adrram[0] ), 
         .Z(n1594)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1461_3_lut.init = 16'hcaca;
    FD1P3AY mem_8__i0_i1 (.D(data[1]), .SP(we_N_63_enable_368), .CK(we_N_63), 
            .Q(\mem[8] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_8__i0_i1.GSR = "ENABLED";
    FD1P3AY mem_7__i0_i7 (.D(data[7]), .SP(we_N_63_enable_377), .CK(we_N_63), 
            .Q(\mem[7] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_7__i0_i7.GSR = "ENABLED";
    FD1P3AY mem_0__i0_i3 (.D(data[3]), .SP(we_N_63_enable_379), .CK(we_N_63), 
            .Q(\mem[0] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_0__i0_i3.GSR = "ENABLED";
    FD1P3AY mem_0__i0_i2 (.D(data[2]), .SP(we_N_63_enable_379), .CK(we_N_63), 
            .Q(\mem[0] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_0__i0_i2.GSR = "ENABLED";
    FD1P3AY mem_7__i0_i6 (.D(data[6]), .SP(we_N_63_enable_377), .CK(we_N_63), 
            .Q(\mem[7] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_7__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_7__i0_i5 (.D(data[5]), .SP(we_N_63_enable_377), .CK(we_N_63), 
            .Q(\mem[7] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_7__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_7__i0_i4 (.D(data[4]), .SP(we_N_63_enable_377), .CK(we_N_63), 
            .Q(\mem[7] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_7__i0_i4.GSR = "ENABLED";
    FD1P3AY mem_7__i0_i3 (.D(data[3]), .SP(we_N_63_enable_377), .CK(we_N_63), 
            .Q(\mem[7] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_7__i0_i3.GSR = "ENABLED";
    FD1P3AY mem_7__i0_i2 (.D(data[2]), .SP(we_N_63_enable_377), .CK(we_N_63), 
            .Q(\mem[7] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_7__i0_i2.GSR = "ENABLED";
    LUT4 i1460_3_lut (.A(\mem[4] [0]), .B(\mem[5] [0]), .C(\adrram[0] ), 
         .Z(n1593)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1460_3_lut.init = 16'hcaca;
    FD1P3AX mem_7__i0_i1 (.D(data[1]), .SP(we_N_63_enable_377), .CK(we_N_63), 
            .Q(\mem[7] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_7__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_6__i0_i7 (.D(data[7]), .SP(we_N_63_enable_386), .CK(we_N_63), 
            .Q(\mem[6] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_6__i0_i7.GSR = "ENABLED";
    FD1P3AY mem_0__i0_i1 (.D(data[1]), .SP(we_N_63_enable_379), .CK(we_N_63), 
            .Q(\mem[0] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_0__i0_i1.GSR = "ENABLED";
    FD1P3AY mem_6__i0_i6 (.D(data[6]), .SP(we_N_63_enable_386), .CK(we_N_63), 
            .Q(\mem[6] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_6__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_6__i0_i5 (.D(data[5]), .SP(we_N_63_enable_386), .CK(we_N_63), 
            .Q(\mem[6] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_6__i0_i5.GSR = "ENABLED";
    FD1P3AY mem_6__i0_i4 (.D(data[4]), .SP(we_N_63_enable_386), .CK(we_N_63), 
            .Q(\mem[6] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_6__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_6__i0_i3 (.D(data[3]), .SP(we_N_63_enable_386), .CK(we_N_63), 
            .Q(\mem[6] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_6__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_63__i0_i7 (.D(data[7]), .SP(we_N_63_enable_405), .CK(we_N_63), 
            .Q(\mem[63] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_63__i0_i7.GSR = "ENABLED";
    LUT4 i1564_3_lut (.A(\mem[26] [3]), .B(\mem[27] [3]), .C(\adrram[0] ), 
         .Z(n1697)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1564_3_lut.init = 16'hcaca;
    FD1P3AX mem_6__i0_i2 (.D(data[2]), .SP(we_N_63_enable_386), .CK(we_N_63), 
            .Q(\mem[6] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_6__i0_i2.GSR = "ENABLED";
    FD1P3AY mem_6__i0_i1 (.D(data[1]), .SP(we_N_63_enable_386), .CK(we_N_63), 
            .Q(\mem[6] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_6__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_63__i0_i6 (.D(data[6]), .SP(we_N_63_enable_405), .CK(we_N_63), 
            .Q(\mem[63] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_63__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_5__i0_i7 (.D(data[7]), .SP(we_N_63_enable_395), .CK(we_N_63), 
            .Q(\mem[5] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_5__i0_i7.GSR = "ENABLED";
    FD1P3AY mem_5__i0_i6 (.D(data[6]), .SP(we_N_63_enable_395), .CK(we_N_63), 
            .Q(\mem[5] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_5__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_5__i0_i5 (.D(data[5]), .SP(we_N_63_enable_395), .CK(we_N_63), 
            .Q(\mem[5] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_5__i0_i5.GSR = "ENABLED";
    FD1P3AY mem_5__i0_i4 (.D(data[4]), .SP(we_N_63_enable_395), .CK(we_N_63), 
            .Q(\mem[5] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_5__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_5__i0_i3 (.D(data[3]), .SP(we_N_63_enable_395), .CK(we_N_63), 
            .Q(\mem[5] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_5__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_63__i0_i5 (.D(data[5]), .SP(we_N_63_enable_405), .CK(we_N_63), 
            .Q(\mem[63] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_63__i0_i5.GSR = "ENABLED";
    LUT4 i1563_3_lut (.A(\mem[24] [3]), .B(\mem[25] [3]), .C(\adrram[0] ), 
         .Z(n1696)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1563_3_lut.init = 16'hcaca;
    FD1P3AY mem_5__i0_i2 (.D(data[2]), .SP(we_N_63_enable_395), .CK(we_N_63), 
            .Q(\mem[5] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_5__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_5__i0_i1 (.D(data[1]), .SP(we_N_63_enable_395), .CK(we_N_63), 
            .Q(\mem[5] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_5__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_63__i0_i4 (.D(data[4]), .SP(we_N_63_enable_405), .CK(we_N_63), 
            .Q(\mem[63] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_63__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_63__i0_i3 (.D(data[3]), .SP(we_N_63_enable_405), .CK(we_N_63), 
            .Q(\mem[63] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_63__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_4__i0_i7 (.D(data[7]), .SP(we_N_63_enable_407), .CK(we_N_63), 
            .Q(\mem[4] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_4__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_4__i0_i6 (.D(data[6]), .SP(we_N_63_enable_407), .CK(we_N_63), 
            .Q(\mem[4] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_4__i0_i6.GSR = "ENABLED";
    FD1P3AY mem_4__i0_i5 (.D(data[5]), .SP(we_N_63_enable_407), .CK(we_N_63), 
            .Q(\mem[4] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_4__i0_i5.GSR = "ENABLED";
    FD1P3AY mem_4__i0_i4 (.D(data[4]), .SP(we_N_63_enable_407), .CK(we_N_63), 
            .Q(\mem[4] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_4__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_63__i0_i2 (.D(data[2]), .SP(we_N_63_enable_405), .CK(we_N_63), 
            .Q(\mem[63] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_63__i0_i2.GSR = "ENABLED";
    LUT4 i1562_3_lut (.A(\mem[22] [3]), .B(\mem[23] [3]), .C(\adrram[0] ), 
         .Z(n1695)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1562_3_lut.init = 16'hcaca;
    FD1P3AY mem_4__i0_i3 (.D(data[3]), .SP(we_N_63_enable_407), .CK(we_N_63), 
            .Q(\mem[4] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_4__i0_i3.GSR = "ENABLED";
    FD1P3AY mem_4__i0_i2 (.D(data[2]), .SP(we_N_63_enable_407), .CK(we_N_63), 
            .Q(\mem[4] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_4__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_63__i0_i1 (.D(data[1]), .SP(we_N_63_enable_405), .CK(we_N_63), 
            .Q(\mem[63] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_63__i0_i1.GSR = "ENABLED";
    FD1P3AY mem_62__i0_i7 (.D(data[7]), .SP(we_N_63_enable_420), .CK(we_N_63), 
            .Q(\mem[62] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_62__i0_i7.GSR = "ENABLED";
    FD1P3AY mem_4__i0_i1 (.D(data[1]), .SP(we_N_63_enable_407), .CK(we_N_63), 
            .Q(\mem[4] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_4__i0_i1.GSR = "ENABLED";
    FD1P3AY mem_3__i0_i7 (.D(data[7]), .SP(we_N_63_enable_416), .CK(we_N_63), 
            .Q(\mem[3] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_3__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_3__i0_i6 (.D(data[6]), .SP(we_N_63_enable_416), .CK(we_N_63), 
            .Q(\mem[3] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_3__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_3__i0_i5 (.D(data[5]), .SP(we_N_63_enable_416), .CK(we_N_63), 
            .Q(\mem[3] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_3__i0_i5.GSR = "ENABLED";
    FD1P3AY mem_62__i0_i6 (.D(data[6]), .SP(we_N_63_enable_420), .CK(we_N_63), 
            .Q(\mem[62] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_62__i0_i6.GSR = "ENABLED";
    LUT4 i1561_3_lut (.A(\mem[20] [3]), .B(\mem[21] [3]), .C(\adrram[0] ), 
         .Z(n1694)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1561_3_lut.init = 16'hcaca;
    FD1P3AY mem_3__i0_i4 (.D(data[4]), .SP(we_N_63_enable_416), .CK(we_N_63), 
            .Q(\mem[3] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_3__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_3__i0_i3 (.D(data[3]), .SP(we_N_63_enable_416), .CK(we_N_63), 
            .Q(\mem[3] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_3__i0_i3.GSR = "ENABLED";
    FD1P3AY mem_62__i0_i5 (.D(data[5]), .SP(we_N_63_enable_420), .CK(we_N_63), 
            .Q(\mem[62] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_62__i0_i5.GSR = "ENABLED";
    FD1P3AY mem_3__i0_i2 (.D(data[2]), .SP(we_N_63_enable_416), .CK(we_N_63), 
            .Q(\mem[3] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_3__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_3__i0_i1 (.D(data[1]), .SP(we_N_63_enable_416), .CK(we_N_63), 
            .Q(\mem[3] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_3__i0_i1.GSR = "ENABLED";
    FD1P3AY mem_62__i0_i4 (.D(data[4]), .SP(we_N_63_enable_420), .CK(we_N_63), 
            .Q(\mem[62] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_62__i0_i4.GSR = "ENABLED";
    LUT4 i1560_3_lut (.A(\mem[18] [3]), .B(\mem[19] [3]), .C(\adrram[0] ), 
         .Z(n1693)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1560_3_lut.init = 16'hcaca;
    LUT4 i1559_3_lut (.A(\mem[16] [3]), .B(\mem[17] [3]), .C(\adrram[0] ), 
         .Z(n1692)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1559_3_lut.init = 16'hcaca;
    LUT4 i1558_3_lut (.A(\mem[14] [3]), .B(\mem[15] [3]), .C(\adrram[0] ), 
         .Z(n1691)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1558_3_lut.init = 16'hcaca;
    FD1P3AY mem_62__i0_i3 (.D(data[3]), .SP(we_N_63_enable_420), .CK(we_N_63), 
            .Q(\mem[62] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_62__i0_i3.GSR = "ENABLED";
    LUT4 i1557_3_lut (.A(\mem[12] [3]), .B(\mem[13] [3]), .C(\adrram[0] ), 
         .Z(n1690)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1557_3_lut.init = 16'hcaca;
    FD1P3AY mem_62__i0_i2 (.D(data[2]), .SP(we_N_63_enable_420), .CK(we_N_63), 
            .Q(\mem[62] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_62__i0_i2.GSR = "ENABLED";
    FD1P3AY mem_62__i0_i1 (.D(data[1]), .SP(we_N_63_enable_420), .CK(we_N_63), 
            .Q(\mem[62] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_62__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_61__i0_i7 (.D(data[7]), .SP(we_N_63_enable_428), .CK(we_N_63), 
            .Q(\mem[61] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_61__i0_i7.GSR = "ENABLED";
    LUT4 i1689_3_lut (.A(\mem[28] [7]), .B(\mem[29] [7]), .C(\adrram[0] ), 
         .Z(n1822)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1689_3_lut.init = 16'hcaca;
    FD1P3AX mem_61__i0_i6 (.D(data[6]), .SP(we_N_63_enable_428), .CK(we_N_63), 
            .Q(\mem[61] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_61__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_61__i0_i5 (.D(data[5]), .SP(we_N_63_enable_428), .CK(we_N_63), 
            .Q(\mem[61] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_61__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_61__i0_i4 (.D(data[4]), .SP(we_N_63_enable_428), .CK(we_N_63), 
            .Q(\mem[61] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_61__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_61__i0_i3 (.D(data[3]), .SP(we_N_63_enable_428), .CK(we_N_63), 
            .Q(\mem[61] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_61__i0_i3.GSR = "ENABLED";
    LUT4 i1932_3_lut (.A(\mem[50] [0]), .B(\mem[51] [0]), .C(\adrram[0] ), 
         .Z(n2065)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1932_3_lut.init = 16'hcaca;
    LUT4 i1814_3_lut (.A(\mem[62] [4]), .B(\mem[63] [4]), .C(\adrram[0] ), 
         .Z(n1947)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1814_3_lut.init = 16'hcaca;
    LUT4 i1934_3_lut (.A(\mem[54] [0]), .B(\mem[55] [0]), .C(\adrram[0] ), 
         .Z(n2067)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1934_3_lut.init = 16'hcaca;
    FD1P3AX mem_61__i0_i2 (.D(data[2]), .SP(we_N_63_enable_428), .CK(we_N_63), 
            .Q(\mem[61] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_61__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_1__i0_i7 (.D(data[7]), .SP(we_N_63_enable_452), .CK(we_N_63), 
            .Q(\mem[1] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_1__i0_i7.GSR = "ENABLED";
    LUT4 i1931_3_lut (.A(\mem[48] [0]), .B(\mem[49] [0]), .C(\adrram[0] ), 
         .Z(n2064)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1931_3_lut.init = 16'hcaca;
    FD1P3AX mem_61__i0_i1 (.D(data[1]), .SP(we_N_63_enable_428), .CK(we_N_63), 
            .Q(\mem[61] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_61__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_60__i0_i7 (.D(data[7]), .SP(we_N_63_enable_437), .CK(we_N_63), 
            .Q(\mem[60] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_60__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_60__i0_i6 (.D(data[6]), .SP(we_N_63_enable_437), .CK(we_N_63), 
            .Q(\mem[60] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_60__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_1__i0_i6 (.D(data[6]), .SP(we_N_63_enable_452), .CK(we_N_63), 
            .Q(\mem[1] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_1__i0_i6.GSR = "ENABLED";
    LUT4 i1813_3_lut (.A(\mem[60] [4]), .B(\mem[61] [4]), .C(\adrram[0] ), 
         .Z(n1946)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1813_3_lut.init = 16'hcaca;
    LUT4 i1803_3_lut (.A(\mem[40] [4]), .B(\mem[41] [4]), .C(\adrram[0] ), 
         .Z(n1936)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1803_3_lut.init = 16'hcaca;
    LUT4 i1933_3_lut (.A(\mem[52] [0]), .B(\mem[53] [0]), .C(\adrram[0] ), 
         .Z(n2066)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1933_3_lut.init = 16'hcaca;
    LUT4 i1930_3_lut (.A(\mem[46] [0]), .B(\mem[47] [0]), .C(\adrram[0] ), 
         .Z(n2063)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1930_3_lut.init = 16'hcaca;
    LUT4 i1926_3_lut (.A(\mem[38] [0]), .B(\mem[39] [0]), .C(\adrram[0] ), 
         .Z(n2059)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1926_3_lut.init = 16'hcaca;
    FD1P3AX mem_60__i0_i5 (.D(data[5]), .SP(we_N_63_enable_437), .CK(we_N_63), 
            .Q(\mem[60] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_60__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_60__i0_i4 (.D(data[4]), .SP(we_N_63_enable_437), .CK(we_N_63), 
            .Q(\mem[60] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_60__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_60__i0_i3 (.D(data[3]), .SP(we_N_63_enable_437), .CK(we_N_63), 
            .Q(\mem[60] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_60__i0_i3.GSR = "ENABLED";
    LUT4 i1688_3_lut (.A(\mem[26] [7]), .B(\mem[27] [7]), .C(\adrram[0] ), 
         .Z(n1821)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1688_3_lut.init = 16'hcaca;
    FD1P3AX mem_60__i0_i2 (.D(data[2]), .SP(we_N_63_enable_437), .CK(we_N_63), 
            .Q(\mem[60] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_60__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_1__i0_i5 (.D(data[5]), .SP(we_N_63_enable_452), .CK(we_N_63), 
            .Q(\mem[1] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_1__i0_i5.GSR = "ENABLED";
    LUT4 i1929_3_lut (.A(\mem[44] [0]), .B(\mem[45] [0]), .C(\adrram[0] ), 
         .Z(n2062)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1929_3_lut.init = 16'hcaca;
    LUT4 i1925_3_lut (.A(\mem[36] [0]), .B(\mem[37] [0]), .C(\adrram[0] ), 
         .Z(n2058)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1925_3_lut.init = 16'hcaca;
    LUT4 i1802_3_lut (.A(\mem[38] [4]), .B(\mem[39] [4]), .C(\adrram[0] ), 
         .Z(n1935)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1802_3_lut.init = 16'hcaca;
    LUT4 i1687_3_lut (.A(\mem[24] [7]), .B(\mem[25] [7]), .C(\adrram[0] ), 
         .Z(n1820)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1687_3_lut.init = 16'hcaca;
    LUT4 i1801_3_lut (.A(\mem[36] [4]), .B(\mem[37] [4]), .C(\adrram[0] ), 
         .Z(n1934)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1801_3_lut.init = 16'hcaca;
    FD1P3AX mem_60__i0_i1 (.D(data[1]), .SP(we_N_63_enable_437), .CK(we_N_63), 
            .Q(\mem[60] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_60__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_59__i0_i7 (.D(data[7]), .SP(we_N_63_enable_446), .CK(we_N_63), 
            .Q(\mem[59] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_59__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_59__i0_i6 (.D(data[6]), .SP(we_N_63_enable_446), .CK(we_N_63), 
            .Q(\mem[59] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_59__i0_i6.GSR = "ENABLED";
    LUT4 i1620_3_lut (.A(\mem[14] [5]), .B(\mem[15] [5]), .C(\adrram[0] ), 
         .Z(n1753)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1620_3_lut.init = 16'hcaca;
    FD1P3AX mem_59__i0_i5 (.D(data[5]), .SP(we_N_63_enable_446), .CK(we_N_63), 
            .Q(\mem[59] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_59__i0_i5.GSR = "ENABLED";
    FD1P3AY mem_1__i0_i4 (.D(data[4]), .SP(we_N_63_enable_452), .CK(we_N_63), 
            .Q(\mem[1] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_1__i0_i4.GSR = "ENABLED";
    LUT4 i1583_3_lut (.A(\mem[2] [4]), .B(\mem[3] [4]), .C(\adrram[0] ), 
         .Z(n1716)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1583_3_lut.init = 16'hcaca;
    LUT4 i1659_3_lut (.A(\mem[30] [6]), .B(\mem[31] [6]), .C(\adrram[0] ), 
         .Z(n1792)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1659_3_lut.init = 16'hcaca;
    LUT4 i1812_3_lut (.A(\mem[58] [4]), .B(\mem[59] [4]), .C(\adrram[0] ), 
         .Z(n1945)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1812_3_lut.init = 16'hcaca;
    LUT4 i1619_3_lut (.A(\mem[12] [5]), .B(\mem[13] [5]), .C(\adrram[0] ), 
         .Z(n1752)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1619_3_lut.init = 16'hcaca;
    LUT4 i2302_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2307), .C(n2314), 
         .D(\adrram[5] ), .Z(we_N_63_enable_336)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2302_2_lut_2_lut_3_lut_4_lut.init = 16'h0002;
    FD1P3AX mem_59__i0_i4 (.D(data[4]), .SP(we_N_63_enable_446), .CK(we_N_63), 
            .Q(\mem[59] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_59__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_59__i0_i3 (.D(data[3]), .SP(we_N_63_enable_446), .CK(we_N_63), 
            .Q(\mem[59] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_59__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_59__i0_i2 (.D(data[2]), .SP(we_N_63_enable_446), .CK(we_N_63), 
            .Q(\mem[59] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_59__i0_i2.GSR = "ENABLED";
    LUT4 i1897_3_lut (.A(\mem[42] [1]), .B(\mem[43] [1]), .C(\adrram[0] ), 
         .Z(n2030)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1897_3_lut.init = 16'hcaca;
    FD1P3AX mem_1__i0_i3 (.D(data[3]), .SP(we_N_63_enable_452), .CK(we_N_63), 
            .Q(\mem[1] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_1__i0_i3.GSR = "ENABLED";
    LUT4 i1658_3_lut (.A(\mem[28] [6]), .B(\mem[29] [6]), .C(\adrram[0] ), 
         .Z(n1791)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1658_3_lut.init = 16'hcaca;
    LUT4 i1811_3_lut (.A(\mem[56] [4]), .B(\mem[57] [4]), .C(\adrram[0] ), 
         .Z(n1944)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1811_3_lut.init = 16'hcaca;
    FD1P3AX mem_59__i0_i1 (.D(data[1]), .SP(we_N_63_enable_446), .CK(we_N_63), 
            .Q(\mem[59] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_59__i0_i1.GSR = "ENABLED";
    LUT4 i1800_3_lut (.A(\mem[34] [4]), .B(\mem[35] [4]), .C(\adrram[0] ), 
         .Z(n1933)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1800_3_lut.init = 16'hcaca;
    LUT4 i1582_3_lut (.A(\mem[0] [4]), .B(\mem[1] [4]), .C(\adrram[0] ), 
         .Z(n1715)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1582_3_lut.init = 16'hcaca;
    FD1P3AX mem_58__i0_i7 (.D(data[7]), .SP(we_N_63_enable_455), .CK(we_N_63), 
            .Q(\mem[58] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_58__i0_i7.GSR = "ENABLED";
    FD1P3AY mem_1__i0_i2 (.D(data[2]), .SP(we_N_63_enable_452), .CK(we_N_63), 
            .Q(\mem[1] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_1__i0_i2.GSR = "ENABLED";
    LUT4 i1502_3_lut (.A(\mem[26] [1]), .B(\mem[27] [1]), .C(\adrram[0] ), 
         .Z(n1635)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1502_3_lut.init = 16'hcaca;
    LUT4 i1896_3_lut (.A(\mem[40] [1]), .B(\mem[41] [1]), .C(\adrram[0] ), 
         .Z(n2029)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1896_3_lut.init = 16'hcaca;
    LUT4 i1799_3_lut (.A(\mem[32] [4]), .B(\mem[33] [4]), .C(\adrram[0] ), 
         .Z(n1932)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1799_3_lut.init = 16'hcaca;
    LUT4 i1618_3_lut (.A(\mem[10] [5]), .B(\mem[11] [5]), .C(\adrram[0] ), 
         .Z(n1751)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1618_3_lut.init = 16'hcaca;
    LUT4 i1501_3_lut (.A(\mem[24] [1]), .B(\mem[25] [1]), .C(\adrram[0] ), 
         .Z(n1634)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1501_3_lut.init = 16'hcaca;
    LUT4 i1928_3_lut (.A(\mem[42] [0]), .B(\mem[43] [0]), .C(\adrram[0] ), 
         .Z(n2061)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1928_3_lut.init = 16'hcaca;
    FD1P3AX mem_58__i0_i6 (.D(data[6]), .SP(we_N_63_enable_455), .CK(we_N_63), 
            .Q(\mem[58] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_58__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_58__i0_i5 (.D(data[5]), .SP(we_N_63_enable_455), .CK(we_N_63), 
            .Q(\mem[58] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_58__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_58__i0_i4 (.D(data[4]), .SP(we_N_63_enable_455), .CK(we_N_63), 
            .Q(\mem[58] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_58__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_1__i0_i1 (.D(data[1]), .SP(we_N_63_enable_452), .CK(we_N_63), 
            .Q(\mem[1] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_1__i0_i1.GSR = "ENABLED";
    LUT4 i1810_3_lut (.A(\mem[54] [4]), .B(\mem[55] [4]), .C(\adrram[0] ), 
         .Z(n1943)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1810_3_lut.init = 16'hcaca;
    FD1P3AX mem_58__i0_i3 (.D(data[3]), .SP(we_N_63_enable_455), .CK(we_N_63), 
            .Q(\mem[58] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_58__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_58__i0_i2 (.D(data[2]), .SP(we_N_63_enable_455), .CK(we_N_63), 
            .Q(\mem[58] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_58__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_58__i0_i1 (.D(data[1]), .SP(we_N_63_enable_455), .CK(we_N_63), 
            .Q(\mem[58] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_58__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_2__i0_i7 (.D(data[7]), .SP(we_N_63_enable_481), .CK(we_N_63), 
            .Q(\mem[2] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_2__i0_i7.GSR = "ENABLED";
    LUT4 i1617_3_lut (.A(\mem[8] [5]), .B(\mem[9] [5]), .C(\adrram[0] ), 
         .Z(n1750)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1617_3_lut.init = 16'hcaca;
    LUT4 i1783_3_lut (.A(\mem[62] [5]), .B(\mem[63] [5]), .C(\adrram[0] ), 
         .Z(n1916)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1783_3_lut.init = 16'hcaca;
    LUT4 i1895_3_lut (.A(\mem[38] [1]), .B(\mem[39] [1]), .C(\adrram[0] ), 
         .Z(n2028)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1895_3_lut.init = 16'hcaca;
    LUT4 i1927_3_lut (.A(\mem[40] [0]), .B(\mem[41] [0]), .C(\adrram[0] ), 
         .Z(n2060)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1927_3_lut.init = 16'hcaca;
    LUT4 i1809_3_lut (.A(\mem[52] [4]), .B(\mem[53] [4]), .C(\adrram[0] ), 
         .Z(n1942)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1809_3_lut.init = 16'hcaca;
    FD1P3AX mem_57__i0_i7 (.D(data[7]), .SP(we_N_63_enable_465), .CK(we_N_63), 
            .Q(\mem[57] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_57__i0_i7.GSR = "ENABLED";
    LUT4 i1628_3_lut (.A(\mem[30] [5]), .B(\mem[31] [5]), .C(\adrram[0] ), 
         .Z(n1761)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1628_3_lut.init = 16'hcaca;
    LUT4 i1782_3_lut (.A(\mem[60] [5]), .B(\mem[61] [5]), .C(\adrram[0] ), 
         .Z(n1915)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1782_3_lut.init = 16'hcaca;
    FD1P3AX mem_57__i0_i6 (.D(data[6]), .SP(we_N_63_enable_465), .CK(we_N_63), 
            .Q(\mem[57] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_57__i0_i6.GSR = "ENABLED";
    FD1P3AY mem_2__i0_i6 (.D(data[6]), .SP(we_N_63_enable_481), .CK(we_N_63), 
            .Q(\mem[2] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_2__i0_i6.GSR = "ENABLED";
    LUT4 i1500_3_lut (.A(\mem[22] [1]), .B(\mem[23] [1]), .C(\adrram[0] ), 
         .Z(n1633)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1500_3_lut.init = 16'hcaca;
    LUT4 i1775_3_lut (.A(\mem[46] [5]), .B(\mem[47] [5]), .C(\adrram[0] ), 
         .Z(n1908)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1775_3_lut.init = 16'hcaca;
    LUT4 i1556_3_lut (.A(\mem[10] [3]), .B(\mem[11] [3]), .C(\adrram[0] ), 
         .Z(n1689)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1556_3_lut.init = 16'hcaca;
    FD1P3AX mem_57__i0_i5 (.D(data[5]), .SP(we_N_63_enable_465), .CK(we_N_63), 
            .Q(\mem[57] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_57__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_57__i0_i4 (.D(data[4]), .SP(we_N_63_enable_465), .CK(we_N_63), 
            .Q(\mem[57] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_57__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_57__i0_i3 (.D(data[3]), .SP(we_N_63_enable_465), .CK(we_N_63), 
            .Q(\mem[57] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_57__i0_i3.GSR = "ENABLED";
    FD1P3AY mem_2__i0_i5 (.D(data[5]), .SP(we_N_63_enable_481), .CK(we_N_63), 
            .Q(\mem[2] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_2__i0_i5.GSR = "ENABLED";
    LUT4 i1894_3_lut (.A(\mem[36] [1]), .B(\mem[37] [1]), .C(\adrram[0] ), 
         .Z(n2027)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1894_3_lut.init = 16'hcaca;
    FD1P3AX mem_57__i0_i2 (.D(data[2]), .SP(we_N_63_enable_465), .CK(we_N_63), 
            .Q(\mem[57] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_57__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_57__i0_i1 (.D(data[1]), .SP(we_N_63_enable_465), .CK(we_N_63), 
            .Q(\mem[57] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_57__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_56__i0_i7 (.D(data[7]), .SP(we_N_63_enable_474), .CK(we_N_63), 
            .Q(\mem[56] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_56__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_56__i0_i6 (.D(data[6]), .SP(we_N_63_enable_474), .CK(we_N_63), 
            .Q(\mem[56] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_56__i0_i6.GSR = "ENABLED";
    FD1P3AY mem_2__i0_i4 (.D(data[4]), .SP(we_N_63_enable_481), .CK(we_N_63), 
            .Q(\mem[2] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_2__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_56__i0_i5 (.D(data[5]), .SP(we_N_63_enable_474), .CK(we_N_63), 
            .Q(\mem[56] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_56__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_56__i0_i4 (.D(data[4]), .SP(we_N_63_enable_474), .CK(we_N_63), 
            .Q(\mem[56] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_56__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_56__i0_i3 (.D(data[3]), .SP(we_N_63_enable_474), .CK(we_N_63), 
            .Q(\mem[56] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_56__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_56__i0_i2 (.D(data[2]), .SP(we_N_63_enable_474), .CK(we_N_63), 
            .Q(\mem[56] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_56__i0_i2.GSR = "ENABLED";
    FD1P3AY mem_2__i0_i3 (.D(data[3]), .SP(we_N_63_enable_481), .CK(we_N_63), 
            .Q(\mem[2] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_2__i0_i3.GSR = "ENABLED";
    LUT4 i1657_3_lut (.A(\mem[26] [6]), .B(\mem[27] [6]), .C(\adrram[0] ), 
         .Z(n1790)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1657_3_lut.init = 16'hcaca;
    FD1P3AX mem_56__i0_i1 (.D(data[1]), .SP(we_N_63_enable_474), .CK(we_N_63), 
            .Q(\mem[56] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_56__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_55__i0_i7 (.D(data[7]), .SP(we_N_63_enable_483), .CK(we_N_63), 
            .Q(\mem[55] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_55__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_55__i0_i6 (.D(data[6]), .SP(we_N_63_enable_483), .CK(we_N_63), 
            .Q(\mem[55] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_55__i0_i6.GSR = "ENABLED";
    FD1P3AY mem_2__i0_i2 (.D(data[2]), .SP(we_N_63_enable_481), .CK(we_N_63), 
            .Q(\mem[2] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_2__i0_i2.GSR = "ENABLED";
    PFUMX i122132_i1 (.BLUT(n1838), .ALUT(n1869), .C0(\adrram[5] ), .Z(data_7__N_66[7]));
    PFUMX i121529_i1 (.BLUT(n1807), .ALUT(n1900), .C0(\adrram[5] ), .Z(data_7__N_66[6]));
    LUT4 i1656_3_lut (.A(\mem[24] [6]), .B(\mem[25] [6]), .C(\adrram[0] ), 
         .Z(n1789)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1656_3_lut.init = 16'hcaca;
    FD1P3AX mem_55__i0_i5 (.D(data[5]), .SP(we_N_63_enable_483), .CK(we_N_63), 
            .Q(\mem[55] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_55__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_55__i0_i4 (.D(data[4]), .SP(we_N_63_enable_483), .CK(we_N_63), 
            .Q(\mem[55] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_55__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_55__i0_i3 (.D(data[3]), .SP(we_N_63_enable_483), .CK(we_N_63), 
            .Q(\mem[55] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_55__i0_i3.GSR = "ENABLED";
    FD1P3AY mem_2__i0_i1 (.D(data[1]), .SP(we_N_63_enable_481), .CK(we_N_63), 
            .Q(\mem[2] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_2__i0_i1.GSR = "ENABLED";
    PFUMX i120926_i1 (.BLUT(n1776), .ALUT(n1931), .C0(\adrram[5] ), .Z(data_7__N_66[5]));
    FD1P3AX mem_55__i0_i2 (.D(data[2]), .SP(we_N_63_enable_483), .CK(we_N_63), 
            .Q(\mem[55] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_55__i0_i2.GSR = "ENABLED";
    PFUMX i120323_i1 (.BLUT(n1745), .ALUT(n1962), .C0(\adrram[5] ), .Z(data_7__N_66[4]));
    FD1P3AX mem_55__i0_i1 (.D(data[1]), .SP(we_N_63_enable_483), .CK(we_N_63), 
            .Q(\mem[55] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_55__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_54__i0_i7 (.D(data[7]), .SP(we_N_63_enable_490), .CK(we_N_63), 
            .Q(\mem[54] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_54__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_54__i0_i6 (.D(data[6]), .SP(we_N_63_enable_490), .CK(we_N_63), 
            .Q(\mem[54] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_54__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_54__i0_i5 (.D(data[5]), .SP(we_N_63_enable_490), .CK(we_N_63), 
            .Q(\mem[54] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_54__i0_i5.GSR = "ENABLED";
    PFUMX i119720_i1 (.BLUT(n1714), .ALUT(n1993), .C0(\adrram[5] ), .Z(data_7__N_66[3]));
    LUT4 i1686_3_lut (.A(\mem[22] [7]), .B(\mem[23] [7]), .C(\adrram[0] ), 
         .Z(n1819)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1686_3_lut.init = 16'hcaca;
    FD1P3AX mem_54__i0_i4 (.D(data[4]), .SP(we_N_63_enable_490), .CK(we_N_63), 
            .Q(\mem[54] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_54__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_54__i0_i3 (.D(data[3]), .SP(we_N_63_enable_490), .CK(we_N_63), 
            .Q(\mem[54] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_54__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_54__i0_i2 (.D(data[2]), .SP(we_N_63_enable_490), .CK(we_N_63), 
            .Q(\mem[54] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_54__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_54__i0_i1 (.D(data[1]), .SP(we_N_63_enable_490), .CK(we_N_63), 
            .Q(\mem[54] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_54__i0_i1.GSR = "ENABLED";
    PFUMX i119117_i1 (.BLUT(n1683), .ALUT(n2024), .C0(\adrram[5] ), .Z(data_7__N_66[2]));
    PFUMX i118514_i1 (.BLUT(n1652), .ALUT(n2055), .C0(\adrram[5] ), .Z(data_7__N_66[1]));
    FD1P3AX mem_53__i0_i7 (.D(data[7]), .SP(we_N_63_enable_497), .CK(we_N_63), 
            .Q(\mem[53] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_53__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_53__i0_i6 (.D(data[6]), .SP(we_N_63_enable_497), .CK(we_N_63), 
            .Q(\mem[53] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_53__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_53__i0_i5 (.D(data[5]), .SP(we_N_63_enable_497), .CK(we_N_63), 
            .Q(\mem[53] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_53__i0_i5.GSR = "ENABLED";
    PFUMX i117911_i1 (.BLUT(n1621), .ALUT(n2086), .C0(\adrram[5] ), .Z(data_7__N_66[0]));
    L6MUX21 i1548 (.D0(n1677), .D1(n1678), .SD(\adrram[3] ), .Z(n1681));
    LUT4 i1685_3_lut (.A(\mem[20] [7]), .B(\mem[21] [7]), .C(\adrram[0] ), 
         .Z(n1818)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1685_3_lut.init = 16'hcaca;
    FD1P3AX mem_53__i0_i4 (.D(data[4]), .SP(we_N_63_enable_497), .CK(we_N_63), 
            .Q(\mem[53] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_53__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_53__i0_i3 (.D(data[3]), .SP(we_N_63_enable_497), .CK(we_N_63), 
            .Q(\mem[53] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_53__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_53__i0_i2 (.D(data[2]), .SP(we_N_63_enable_497), .CK(we_N_63), 
            .Q(\mem[53] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_53__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_53__i0_i1 (.D(data[1]), .SP(we_N_63_enable_497), .CK(we_N_63), 
            .Q(\mem[53] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_53__i0_i1.GSR = "ENABLED";
    L6MUX21 i1549 (.D0(n1679), .D1(n1680), .SD(\adrram[3] ), .Z(n1682));
    L6MUX21 i1486 (.D0(n1615), .D1(n1616), .SD(\adrram[3] ), .Z(n1619));
    L6MUX21 i1611 (.D0(n1741), .D1(n1742), .SD(\adrram[3] ), .Z(n1744));
    L6MUX21 i1610 (.D0(n1739), .D1(n1740), .SD(\adrram[3] ), .Z(n1743));
    L6MUX21 i1734 (.D0(n1863), .D1(n1864), .SD(\adrram[3] ), .Z(n1867));
    LUT4 i1808_3_lut (.A(\mem[50] [4]), .B(\mem[51] [4]), .C(\adrram[0] ), 
         .Z(n1941)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1808_3_lut.init = 16'hcaca;
    FD1P3AX mem_52__i0_i7 (.D(data[7]), .SP(we_N_63_enable_504), .CK(we_N_63), 
            .Q(\mem[52] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_52__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_52__i0_i6 (.D(data[6]), .SP(we_N_63_enable_504), .CK(we_N_63), 
            .Q(\mem[52] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_52__i0_i6.GSR = "ENABLED";
    FD1P3AX mem_52__i0_i5 (.D(data[5]), .SP(we_N_63_enable_504), .CK(we_N_63), 
            .Q(\mem[52] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_52__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_52__i0_i4 (.D(data[4]), .SP(we_N_63_enable_504), .CK(we_N_63), 
            .Q(\mem[52] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_52__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_52__i0_i3 (.D(data[3]), .SP(we_N_63_enable_504), .CK(we_N_63), 
            .Q(\mem[52] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_52__i0_i3.GSR = "ENABLED";
    L6MUX21 i1735 (.D0(n1865), .D1(n1866), .SD(\adrram[3] ), .Z(n1868));
    L6MUX21 i1858 (.D0(n1987), .D1(n1988), .SD(\adrram[3] ), .Z(n1991));
    L6MUX21 i1859 (.D0(n1989), .D1(n1990), .SD(\adrram[3] ), .Z(n1992));
    L6MUX21 i1920 (.D0(n2049), .D1(n2050), .SD(\adrram[3] ), .Z(n2053));
    LUT4 i1627_3_lut (.A(\mem[28] [5]), .B(\mem[29] [5]), .C(\adrram[0] ), 
         .Z(n1760)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1627_3_lut.init = 16'hcaca;
    FD1P3AX mem_52__i0_i2 (.D(data[2]), .SP(we_N_63_enable_504), .CK(we_N_63), 
            .Q(\mem[52] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_52__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_52__i0_i1 (.D(data[1]), .SP(we_N_63_enable_504), .CK(we_N_63), 
            .Q(\mem[52] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_52__i0_i1.GSR = "ENABLED";
    FD1P3AX mem_51__i0_i7 (.D(data[7]), .SP(we_N_63_enable_511), .CK(we_N_63), 
            .Q(\mem[51] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_51__i0_i7.GSR = "ENABLED";
    FD1P3AX mem_51__i0_i6 (.D(data[6]), .SP(we_N_63_enable_511), .CK(we_N_63), 
            .Q(\mem[51] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_51__i0_i6.GSR = "ENABLED";
    L6MUX21 i1921 (.D0(n2051), .D1(n2052), .SD(\adrram[3] ), .Z(n2054));
    L6MUX21 i1951 (.D0(n2080), .D1(n2081), .SD(\adrram[3] ), .Z(n2084));
    L6MUX21 i1952 (.D0(n2082), .D1(n2083), .SD(\adrram[3] ), .Z(n2085));
    L6MUX21 i1765 (.D0(n1894), .D1(n1895), .SD(\adrram[3] ), .Z(n1898));
    LUT4 i1655_3_lut (.A(\mem[22] [6]), .B(\mem[23] [6]), .C(\adrram[0] ), 
         .Z(n1788)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1655_3_lut.init = 16'hcaca;
    FD1P3AX mem_51__i0_i5 (.D(data[5]), .SP(we_N_63_enable_511), .CK(we_N_63), 
            .Q(\mem[51] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_51__i0_i5.GSR = "ENABLED";
    FD1P3AX mem_51__i0_i4 (.D(data[4]), .SP(we_N_63_enable_511), .CK(we_N_63), 
            .Q(\mem[51] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_51__i0_i4.GSR = "ENABLED";
    FD1P3AX mem_51__i0_i3 (.D(data[3]), .SP(we_N_63_enable_511), .CK(we_N_63), 
            .Q(\mem[51] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_51__i0_i3.GSR = "ENABLED";
    FD1P3AX mem_51__i0_i2 (.D(data[2]), .SP(we_N_63_enable_511), .CK(we_N_63), 
            .Q(\mem[51] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_51__i0_i2.GSR = "ENABLED";
    FD1P3AX mem_51__i0_i1 (.D(data[1]), .SP(we_N_63_enable_511), .CK(we_N_63), 
            .Q(\mem[51] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_51__i0_i1.GSR = "ENABLED";
    L6MUX21 i1766 (.D0(n1896), .D1(n1897), .SD(\adrram[3] ), .Z(n1899));
    L6MUX21 i1517 (.D0(n1646), .D1(n1647), .SD(\adrram[3] ), .Z(n1650));
    L6MUX21 i1518 (.D0(n1648), .D1(n1649), .SD(\adrram[3] ), .Z(n1651));
    L6MUX21 i1487 (.D0(n1617), .D1(n1618), .SD(\adrram[3] ), .Z(n1620));
    LUT4 i1684_3_lut (.A(\mem[18] [7]), .B(\mem[19] [7]), .C(\adrram[0] ), 
         .Z(n1817)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1684_3_lut.init = 16'hcaca;
    L6MUX21 i1579 (.D0(n1708), .D1(n1709), .SD(\adrram[3] ), .Z(n1712));
    LUT4 i1654_3_lut (.A(\mem[20] [6]), .B(\mem[21] [6]), .C(\adrram[0] ), 
         .Z(n1787)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1654_3_lut.init = 16'hcaca;
    PFUMX i1945 (.BLUT(n2068), .ALUT(n2069), .C0(\adrram[1] ), .Z(n2078));
    PFUMX i1512 (.BLUT(n1636), .ALUT(n1637), .C0(\adrram[1] ), .Z(n1645));
    LUT4 i1807_3_lut (.A(\mem[48] [4]), .B(\mem[49] [4]), .C(\adrram[0] ), 
         .Z(n1940)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1807_3_lut.init = 16'hcaca;
    LUT4 i1683_3_lut (.A(\mem[16] [7]), .B(\mem[17] [7]), .C(\adrram[0] ), 
         .Z(n1816)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1683_3_lut.init = 16'hcaca;
    LUT4 i1653_3_lut (.A(\mem[18] [6]), .B(\mem[19] [6]), .C(\adrram[0] ), 
         .Z(n1786)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1653_3_lut.init = 16'hcaca;
    LUT4 i1616_3_lut (.A(\mem[6] [5]), .B(\mem[7] [5]), .C(\adrram[0] ), 
         .Z(n1749)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1616_3_lut.init = 16'hcaca;
    LUT4 i1652_3_lut (.A(\mem[16] [6]), .B(\mem[17] [6]), .C(\adrram[0] ), 
         .Z(n1785)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1652_3_lut.init = 16'hcaca;
    LUT4 i1682_3_lut (.A(\mem[14] [7]), .B(\mem[15] [7]), .C(\adrram[0] ), 
         .Z(n1815)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1682_3_lut.init = 16'hcaca;
    LUT4 i1681_3_lut (.A(\mem[12] [7]), .B(\mem[13] [7]), .C(\adrram[0] ), 
         .Z(n1814)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1681_3_lut.init = 16'hcaca;
    LUT4 i1806_3_lut (.A(\mem[46] [4]), .B(\mem[47] [4]), .C(\adrram[0] ), 
         .Z(n1939)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1806_3_lut.init = 16'hcaca;
    LUT4 i1626_3_lut (.A(\mem[26] [5]), .B(\mem[27] [5]), .C(\adrram[0] ), 
         .Z(n1759)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1626_3_lut.init = 16'hcaca;
    LUT4 i1651_3_lut (.A(\mem[14] [6]), .B(\mem[15] [6]), .C(\adrram[0] ), 
         .Z(n1784)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1651_3_lut.init = 16'hcaca;
    LUT4 i1680_3_lut (.A(\mem[10] [7]), .B(\mem[11] [7]), .C(\adrram[0] ), 
         .Z(n1813)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1680_3_lut.init = 16'hcaca;
    LUT4 i1650_3_lut (.A(\mem[12] [6]), .B(\mem[13] [6]), .C(\adrram[0] ), 
         .Z(n1783)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1650_3_lut.init = 16'hcaca;
    LUT4 i1805_3_lut (.A(\mem[44] [4]), .B(\mem[45] [4]), .C(\adrram[0] ), 
         .Z(n1938)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1805_3_lut.init = 16'hcaca;
    LUT4 i1625_3_lut (.A(\mem[24] [5]), .B(\mem[25] [5]), .C(\adrram[0] ), 
         .Z(n1758)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1625_3_lut.init = 16'hcaca;
    LUT4 i1615_3_lut (.A(\mem[4] [5]), .B(\mem[5] [5]), .C(\adrram[0] ), 
         .Z(n1748)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1615_3_lut.init = 16'hcaca;
    LUT4 i1679_3_lut (.A(\mem[8] [7]), .B(\mem[9] [7]), .C(\adrram[0] ), 
         .Z(n1812)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1679_3_lut.init = 16'hcaca;
    LUT4 i1649_3_lut (.A(\mem[10] [6]), .B(\mem[11] [6]), .C(\adrram[0] ), 
         .Z(n1782)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1649_3_lut.init = 16'hcaca;
    LUT4 i1648_3_lut (.A(\mem[8] [6]), .B(\mem[9] [6]), .C(\adrram[0] ), 
         .Z(n1781)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1648_3_lut.init = 16'hcaca;
    LUT4 i1678_3_lut (.A(\mem[6] [7]), .B(\mem[7] [7]), .C(\adrram[0] ), 
         .Z(n1811)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1678_3_lut.init = 16'hcaca;
    LUT4 i1677_3_lut (.A(\mem[4] [7]), .B(\mem[5] [7]), .C(\adrram[0] ), 
         .Z(n1810)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1677_3_lut.init = 16'hcaca;
    LUT4 i1924_3_lut (.A(\mem[34] [0]), .B(\mem[35] [0]), .C(\adrram[0] ), 
         .Z(n2057)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1924_3_lut.init = 16'hcaca;
    PFUMX i1846 (.BLUT(n1963), .ALUT(n1964), .C0(\adrram[1] ), .Z(n1979));
    LUT4 i1624_3_lut (.A(\mem[22] [5]), .B(\mem[23] [5]), .C(\adrram[0] ), 
         .Z(n1757)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1624_3_lut.init = 16'hcaca;
    LUT4 i1614_3_lut (.A(\mem[2] [5]), .B(\mem[3] [5]), .C(\adrram[0] ), 
         .Z(n1747)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1614_3_lut.init = 16'hcaca;
    LUT4 i1471_3_lut (.A(\mem[26] [0]), .B(\mem[27] [0]), .C(\adrram[0] ), 
         .Z(n1604)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1471_3_lut.init = 16'hcaca;
    LUT4 i1499_3_lut (.A(\mem[20] [1]), .B(\mem[21] [1]), .C(\adrram[0] ), 
         .Z(n1632)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1499_3_lut.init = 16'hcaca;
    LUT4 i1647_3_lut (.A(\mem[6] [6]), .B(\mem[7] [6]), .C(\adrram[0] ), 
         .Z(n1780)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1647_3_lut.init = 16'hcaca;
    LUT4 i1676_3_lut (.A(\mem[2] [7]), .B(\mem[3] [7]), .C(\adrram[0] ), 
         .Z(n1809)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1676_3_lut.init = 16'hcaca;
    LUT4 i1646_3_lut (.A(\mem[4] [6]), .B(\mem[5] [6]), .C(\adrram[0] ), 
         .Z(n1779)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1646_3_lut.init = 16'hcaca;
    LUT4 i1923_3_lut (.A(\mem[32] [0]), .B(\mem[33] [0]), .C(\adrram[0] ), 
         .Z(n2056)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1923_3_lut.init = 16'hcaca;
    LUT4 i1623_3_lut (.A(\mem[20] [5]), .B(\mem[21] [5]), .C(\adrram[0] ), 
         .Z(n1756)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1623_3_lut.init = 16'hcaca;
    LUT4 i1613_3_lut (.A(\mem[0] [5]), .B(\mem[1] [5]), .C(\adrram[0] ), 
         .Z(n1746)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1613_3_lut.init = 16'hcaca;
    LUT4 i1470_3_lut (.A(\mem[24] [0]), .B(\mem[25] [0]), .C(\adrram[0] ), 
         .Z(n1603)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1470_3_lut.init = 16'hcaca;
    LUT4 i1774_3_lut (.A(\mem[44] [5]), .B(\mem[45] [5]), .C(\adrram[0] ), 
         .Z(n1907)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1774_3_lut.init = 16'hcaca;
    LUT4 i1675_3_lut (.A(\mem[0] [7]), .B(\mem[1] [7]), .C(\adrram[0] ), 
         .Z(n1808)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1675_3_lut.init = 16'hcaca;
    LUT4 i1645_3_lut (.A(\mem[2] [6]), .B(\mem[3] [6]), .C(\adrram[0] ), 
         .Z(n1778)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1645_3_lut.init = 16'hcaca;
    LUT4 i1779_3_lut (.A(\mem[54] [5]), .B(\mem[55] [5]), .C(\adrram[0] ), 
         .Z(n1912)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1779_3_lut.init = 16'hcaca;
    LUT4 i1644_3_lut (.A(\mem[0] [6]), .B(\mem[1] [6]), .C(\adrram[0] ), 
         .Z(n1777)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1644_3_lut.init = 16'hcaca;
    LUT4 i1893_3_lut (.A(\mem[34] [1]), .B(\mem[35] [1]), .C(\adrram[0] ), 
         .Z(n2026)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1893_3_lut.init = 16'hcaca;
    LUT4 i1892_3_lut (.A(\mem[32] [1]), .B(\mem[33] [1]), .C(\adrram[0] ), 
         .Z(n2025)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1892_3_lut.init = 16'hcaca;
    LUT4 i1804_3_lut (.A(\mem[42] [4]), .B(\mem[43] [4]), .C(\adrram[0] ), 
         .Z(n1937)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1804_3_lut.init = 16'hcaca;
    LUT4 i1622_3_lut (.A(\mem[18] [5]), .B(\mem[19] [5]), .C(\adrram[0] ), 
         .Z(n1755)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1622_3_lut.init = 16'hcaca;
    LUT4 i1585_3_lut (.A(\mem[6] [4]), .B(\mem[7] [4]), .C(\adrram[0] ), 
         .Z(n1718)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1585_3_lut.init = 16'hcaca;
    LUT4 i1781_3_lut (.A(\mem[58] [5]), .B(\mem[59] [5]), .C(\adrram[0] ), 
         .Z(n1914)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1781_3_lut.init = 16'hcaca;
    LUT4 i1778_3_lut (.A(\mem[52] [5]), .B(\mem[53] [5]), .C(\adrram[0] ), 
         .Z(n1911)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1778_3_lut.init = 16'hcaca;
    LUT4 i1555_3_lut (.A(\mem[8] [3]), .B(\mem[9] [3]), .C(\adrram[0] ), 
         .Z(n1688)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1555_3_lut.init = 16'hcaca;
    LUT4 i1714_3_lut (.A(\mem[48] [7]), .B(\mem[49] [7]), .C(\adrram[0] ), 
         .Z(n1847)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1714_3_lut.init = 16'hcaca;
    LUT4 i1715_3_lut (.A(\mem[50] [7]), .B(\mem[51] [7]), .C(\adrram[0] ), 
         .Z(n1848)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1715_3_lut.init = 16'hcaca;
    LUT4 i1844_3_lut (.A(\mem[60] [3]), .B(\mem[61] [3]), .C(\adrram[0] ), 
         .Z(n1977)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1844_3_lut.init = 16'hcaca;
    LUT4 i1845_3_lut (.A(\mem[62] [3]), .B(\mem[63] [3]), .C(\adrram[0] ), 
         .Z(n1978)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1845_3_lut.init = 16'hcaca;
    LUT4 i1716_3_lut (.A(\mem[52] [7]), .B(\mem[53] [7]), .C(\adrram[0] ), 
         .Z(n1849)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1716_3_lut.init = 16'hcaca;
    LUT4 i1717_3_lut (.A(\mem[54] [7]), .B(\mem[55] [7]), .C(\adrram[0] ), 
         .Z(n1850)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1717_3_lut.init = 16'hcaca;
    LUT4 i1718_3_lut (.A(\mem[56] [7]), .B(\mem[57] [7]), .C(\adrram[0] ), 
         .Z(n1851)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1718_3_lut.init = 16'hcaca;
    LUT4 i1719_3_lut (.A(\mem[58] [7]), .B(\mem[59] [7]), .C(\adrram[0] ), 
         .Z(n1852)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1719_3_lut.init = 16'hcaca;
    LUT4 i1720_3_lut (.A(\mem[60] [7]), .B(\mem[61] [7]), .C(\adrram[0] ), 
         .Z(n1853)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1720_3_lut.init = 16'hcaca;
    LUT4 i1721_3_lut (.A(\mem[62] [7]), .B(\mem[63] [7]), .C(\adrram[0] ), 
         .Z(n1854)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1721_3_lut.init = 16'hcaca;
    LUT4 i1596_3_lut (.A(\mem[28] [4]), .B(\mem[29] [4]), .C(\adrram[0] ), 
         .Z(n1729)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1596_3_lut.init = 16'hcaca;
    LUT4 i1597_3_lut (.A(\mem[30] [4]), .B(\mem[31] [4]), .C(\adrram[0] ), 
         .Z(n1730)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1597_3_lut.init = 16'hcaca;
    LUT4 i1594_3_lut (.A(\mem[24] [4]), .B(\mem[25] [4]), .C(\adrram[0] ), 
         .Z(n1727)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1594_3_lut.init = 16'hcaca;
    LUT4 i1595_3_lut (.A(\mem[26] [4]), .B(\mem[27] [4]), .C(\adrram[0] ), 
         .Z(n1728)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1595_3_lut.init = 16'hcaca;
    LUT4 i1592_3_lut (.A(\mem[20] [4]), .B(\mem[21] [4]), .C(\adrram[0] ), 
         .Z(n1725)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1592_3_lut.init = 16'hcaca;
    LUT4 i1593_3_lut (.A(\mem[22] [4]), .B(\mem[23] [4]), .C(\adrram[0] ), 
         .Z(n1726)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1593_3_lut.init = 16'hcaca;
    LUT4 i1590_3_lut (.A(\mem[16] [4]), .B(\mem[17] [4]), .C(\adrram[0] ), 
         .Z(n1723)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1590_3_lut.init = 16'hcaca;
    LUT4 i1591_3_lut (.A(\mem[18] [4]), .B(\mem[19] [4]), .C(\adrram[0] ), 
         .Z(n1724)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1591_3_lut.init = 16'hcaca;
    LUT4 i1588_3_lut (.A(\mem[12] [4]), .B(\mem[13] [4]), .C(\adrram[0] ), 
         .Z(n1721)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1588_3_lut.init = 16'hcaca;
    LUT4 i1589_3_lut (.A(\mem[14] [4]), .B(\mem[15] [4]), .C(\adrram[0] ), 
         .Z(n1722)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1589_3_lut.init = 16'hcaca;
    LUT4 i1586_3_lut (.A(\mem[8] [4]), .B(\mem[9] [4]), .C(\adrram[0] ), 
         .Z(n1719)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1586_3_lut.init = 16'hcaca;
    LUT4 i1587_3_lut (.A(\mem[10] [4]), .B(\mem[11] [4]), .C(\adrram[0] ), 
         .Z(n1720)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1587_3_lut.init = 16'hcaca;
    LUT4 i1458_3_lut (.A(\mem[0] [0]), .B(\mem[1] [0]), .C(\adrram[0] ), 
         .Z(n1591)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1458_3_lut.init = 16'hcaca;
    LUT4 i1459_3_lut (.A(\mem[2] [0]), .B(\mem[3] [0]), .C(\adrram[0] ), 
         .Z(n1592)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1459_3_lut.init = 16'hcaca;
    LUT4 i1621_3_lut (.A(\mem[16] [5]), .B(\mem[17] [5]), .C(\adrram[0] ), 
         .Z(n1754)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1621_3_lut.init = 16'hcaca;
    LUT4 i1584_3_lut (.A(\mem[4] [4]), .B(\mem[5] [4]), .C(\adrram[0] ), 
         .Z(n1717)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1584_3_lut.init = 16'hcaca;
    LUT4 i1874_3_lut (.A(\mem[58] [2]), .B(\mem[59] [2]), .C(\adrram[0] ), 
         .Z(n2007)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1874_3_lut.init = 16'hcaca;
    LUT4 i1876_3_lut (.A(\mem[62] [2]), .B(\mem[63] [2]), .C(\adrram[0] ), 
         .Z(n2009)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1876_3_lut.init = 16'hcaca;
    LUT4 i1875_3_lut (.A(\mem[60] [2]), .B(\mem[61] [2]), .C(\adrram[0] ), 
         .Z(n2008)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1875_3_lut.init = 16'hcaca;
    LUT4 i1498_3_lut (.A(\mem[18] [1]), .B(\mem[19] [1]), .C(\adrram[0] ), 
         .Z(n1631)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1498_3_lut.init = 16'hcaca;
    LUT4 i1497_3_lut (.A(\mem[16] [1]), .B(\mem[17] [1]), .C(\adrram[0] ), 
         .Z(n1630)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1497_3_lut.init = 16'hcaca;
    LUT4 i1554_3_lut (.A(\mem[6] [3]), .B(\mem[7] [3]), .C(\adrram[0] ), 
         .Z(n1687)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1554_3_lut.init = 16'hcaca;
    LUT4 i1553_3_lut (.A(\mem[4] [3]), .B(\mem[5] [3]), .C(\adrram[0] ), 
         .Z(n1686)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1553_3_lut.init = 16'hcaca;
    LUT4 i1552_3_lut (.A(\mem[2] [3]), .B(\mem[3] [3]), .C(\adrram[0] ), 
         .Z(n1685)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1552_3_lut.init = 16'hcaca;
    LUT4 i1551_3_lut (.A(\mem[0] [3]), .B(\mem[1] [3]), .C(\adrram[0] ), 
         .Z(n1684)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1551_3_lut.init = 16'hcaca;
    LUT4 i1752_3_lut (.A(\mem[62] [6]), .B(\mem[63] [6]), .C(\adrram[0] ), 
         .Z(n1885)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1752_3_lut.init = 16'hcaca;
    LUT4 i1751_3_lut (.A(\mem[60] [6]), .B(\mem[61] [6]), .C(\adrram[0] ), 
         .Z(n1884)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1751_3_lut.init = 16'hcaca;
    LUT4 i1750_3_lut (.A(\mem[58] [6]), .B(\mem[59] [6]), .C(\adrram[0] ), 
         .Z(n1883)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1750_3_lut.init = 16'hcaca;
    LUT4 i1749_3_lut (.A(\mem[56] [6]), .B(\mem[57] [6]), .C(\adrram[0] ), 
         .Z(n1882)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1749_3_lut.init = 16'hcaca;
    LUT4 i1748_3_lut (.A(\mem[54] [6]), .B(\mem[55] [6]), .C(\adrram[0] ), 
         .Z(n1881)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1748_3_lut.init = 16'hcaca;
    LUT4 i1747_3_lut (.A(\mem[52] [6]), .B(\mem[53] [6]), .C(\adrram[0] ), 
         .Z(n1880)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1747_3_lut.init = 16'hcaca;
    LUT4 i1777_3_lut (.A(\mem[50] [5]), .B(\mem[51] [5]), .C(\adrram[0] ), 
         .Z(n1910)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1777_3_lut.init = 16'hcaca;
    LUT4 i1776_3_lut (.A(\mem[48] [5]), .B(\mem[49] [5]), .C(\adrram[0] ), 
         .Z(n1909)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1776_3_lut.init = 16'hcaca;
    LUT4 i1873_3_lut (.A(\mem[56] [2]), .B(\mem[57] [2]), .C(\adrram[0] ), 
         .Z(n2006)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1873_3_lut.init = 16'hcaca;
    LUT4 i1496_3_lut (.A(\mem[14] [1]), .B(\mem[15] [1]), .C(\adrram[0] ), 
         .Z(n1629)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1496_3_lut.init = 16'hcaca;
    LUT4 i1495_3_lut (.A(\mem[12] [1]), .B(\mem[13] [1]), .C(\adrram[0] ), 
         .Z(n1628)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1495_3_lut.init = 16'hcaca;
    LUT4 i1492_3_lut (.A(\mem[6] [1]), .B(\mem[7] [1]), .C(\adrram[0] ), 
         .Z(n1625)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1492_3_lut.init = 16'hcaca;
    LUT4 i1491_3_lut (.A(\mem[4] [1]), .B(\mem[5] [1]), .C(\adrram[0] ), 
         .Z(n1624)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1491_3_lut.init = 16'hcaca;
    LUT4 i1490_3_lut (.A(\mem[2] [1]), .B(\mem[3] [1]), .C(\adrram[0] ), 
         .Z(n1623)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1490_3_lut.init = 16'hcaca;
    LUT4 i1780_3_lut (.A(\mem[56] [5]), .B(\mem[57] [5]), .C(\adrram[0] ), 
         .Z(n1913)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1780_3_lut.init = 16'hcaca;
    LUT4 i1494_3_lut (.A(\mem[10] [1]), .B(\mem[11] [1]), .C(\adrram[0] ), 
         .Z(n1627)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1494_3_lut.init = 16'hcaca;
    LUT4 i1489_3_lut (.A(\mem[0] [1]), .B(\mem[1] [1]), .C(\adrram[0] ), 
         .Z(n1622)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1489_3_lut.init = 16'hcaca;
    LUT4 i1493_3_lut (.A(\mem[8] [1]), .B(\mem[9] [1]), .C(\adrram[0] ), 
         .Z(n1626)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1493_3_lut.init = 16'hcaca;
    LUT4 i1773_3_lut (.A(\mem[42] [5]), .B(\mem[43] [5]), .C(\adrram[0] ), 
         .Z(n1906)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1773_3_lut.init = 16'hcaca;
    LUT4 i1772_3_lut (.A(\mem[40] [5]), .B(\mem[41] [5]), .C(\adrram[0] ), 
         .Z(n1905)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1772_3_lut.init = 16'hcaca;
    LUT4 i1746_3_lut (.A(\mem[50] [6]), .B(\mem[51] [6]), .C(\adrram[0] ), 
         .Z(n1879)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1746_3_lut.init = 16'hcaca;
    LUT4 i1745_3_lut (.A(\mem[48] [6]), .B(\mem[49] [6]), .C(\adrram[0] ), 
         .Z(n1878)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1745_3_lut.init = 16'hcaca;
    LUT4 i1744_3_lut (.A(\mem[46] [6]), .B(\mem[47] [6]), .C(\adrram[0] ), 
         .Z(n1877)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1744_3_lut.init = 16'hcaca;
    LUT4 i1743_3_lut (.A(\mem[44] [6]), .B(\mem[45] [6]), .C(\adrram[0] ), 
         .Z(n1876)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1743_3_lut.init = 16'hcaca;
    LUT4 i1742_3_lut (.A(\mem[42] [6]), .B(\mem[43] [6]), .C(\adrram[0] ), 
         .Z(n1875)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1742_3_lut.init = 16'hcaca;
    LUT4 i1741_3_lut (.A(\mem[40] [6]), .B(\mem[41] [6]), .C(\adrram[0] ), 
         .Z(n1874)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1741_3_lut.init = 16'hcaca;
    LUT4 i1740_3_lut (.A(\mem[38] [6]), .B(\mem[39] [6]), .C(\adrram[0] ), 
         .Z(n1873)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1740_3_lut.init = 16'hcaca;
    LUT4 i1739_3_lut (.A(\mem[36] [6]), .B(\mem[37] [6]), .C(\adrram[0] ), 
         .Z(n1872)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1739_3_lut.init = 16'hcaca;
    LUT4 i1738_3_lut (.A(\mem[34] [6]), .B(\mem[35] [6]), .C(\adrram[0] ), 
         .Z(n1871)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1738_3_lut.init = 16'hcaca;
    LUT4 i1737_3_lut (.A(\mem[32] [6]), .B(\mem[33] [6]), .C(\adrram[0] ), 
         .Z(n1870)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1737_3_lut.init = 16'hcaca;
    LUT4 i1713_3_lut (.A(\mem[46] [7]), .B(\mem[47] [7]), .C(\adrram[0] ), 
         .Z(n1846)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1713_3_lut.init = 16'hcaca;
    PFUMX i1911 (.BLUT(n2031), .ALUT(n2032), .C0(\adrram[1] ), .Z(n2044));
    LUT4 i1712_3_lut (.A(\mem[44] [7]), .B(\mem[45] [7]), .C(\adrram[0] ), 
         .Z(n1845)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1712_3_lut.init = 16'hcaca;
    LUT4 i1843_3_lut (.A(\mem[58] [3]), .B(\mem[59] [3]), .C(\adrram[0] ), 
         .Z(n1976)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1843_3_lut.init = 16'hcaca;
    LUT4 i1842_3_lut (.A(\mem[56] [3]), .B(\mem[57] [3]), .C(\adrram[0] ), 
         .Z(n1975)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1842_3_lut.init = 16'hcaca;
    LUT4 i1711_3_lut (.A(\mem[42] [7]), .B(\mem[43] [7]), .C(\adrram[0] ), 
         .Z(n1844)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1711_3_lut.init = 16'hcaca;
    LUT4 i1710_3_lut (.A(\mem[40] [7]), .B(\mem[41] [7]), .C(\adrram[0] ), 
         .Z(n1843)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1710_3_lut.init = 16'hcaca;
    LUT4 i1709_3_lut (.A(\mem[38] [7]), .B(\mem[39] [7]), .C(\adrram[0] ), 
         .Z(n1842)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1709_3_lut.init = 16'hcaca;
    LUT4 i1708_3_lut (.A(\mem[36] [7]), .B(\mem[37] [7]), .C(\adrram[0] ), 
         .Z(n1841)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1708_3_lut.init = 16'hcaca;
    LUT4 i1841_3_lut (.A(\mem[54] [3]), .B(\mem[55] [3]), .C(\adrram[0] ), 
         .Z(n1974)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1841_3_lut.init = 16'hcaca;
    LUT4 i1840_3_lut (.A(\mem[52] [3]), .B(\mem[53] [3]), .C(\adrram[0] ), 
         .Z(n1973)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1840_3_lut.init = 16'hcaca;
    LUT4 i1907_3_lut (.A(\mem[62] [1]), .B(\mem[63] [1]), .C(\adrram[0] ), 
         .Z(n2040)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1907_3_lut.init = 16'hcaca;
    LUT4 i1906_3_lut (.A(\mem[60] [1]), .B(\mem[61] [1]), .C(\adrram[0] ), 
         .Z(n2039)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1906_3_lut.init = 16'hcaca;
    LUT4 i1707_3_lut (.A(\mem[34] [7]), .B(\mem[35] [7]), .C(\adrram[0] ), 
         .Z(n1840)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1707_3_lut.init = 16'hcaca;
    LUT4 i1706_3_lut (.A(\mem[32] [7]), .B(\mem[33] [7]), .C(\adrram[0] ), 
         .Z(n1839)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1706_3_lut.init = 16'hcaca;
    LUT4 i1839_3_lut (.A(\mem[50] [3]), .B(\mem[51] [3]), .C(\adrram[0] ), 
         .Z(n1972)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1839_3_lut.init = 16'hcaca;
    LUT4 i1838_3_lut (.A(\mem[48] [3]), .B(\mem[49] [3]), .C(\adrram[0] ), 
         .Z(n1971)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1838_3_lut.init = 16'hcaca;
    LUT4 i1837_3_lut (.A(\mem[46] [3]), .B(\mem[47] [3]), .C(\adrram[0] ), 
         .Z(n1970)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1837_3_lut.init = 16'hcaca;
    LUT4 i1836_3_lut (.A(\mem[44] [3]), .B(\mem[45] [3]), .C(\adrram[0] ), 
         .Z(n1969)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1836_3_lut.init = 16'hcaca;
    LUT4 i1905_3_lut (.A(\mem[58] [1]), .B(\mem[59] [1]), .C(\adrram[0] ), 
         .Z(n2038)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1905_3_lut.init = 16'hcaca;
    LUT4 i1904_3_lut (.A(\mem[56] [1]), .B(\mem[57] [1]), .C(\adrram[0] ), 
         .Z(n2037)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1904_3_lut.init = 16'hcaca;
    LUT4 i1835_3_lut (.A(\mem[42] [3]), .B(\mem[43] [3]), .C(\adrram[0] ), 
         .Z(n1968)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1835_3_lut.init = 16'hcaca;
    LUT4 i1834_3_lut (.A(\mem[40] [3]), .B(\mem[41] [3]), .C(\adrram[0] ), 
         .Z(n1967)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1834_3_lut.init = 16'hcaca;
    LUT4 i1535_3_lut (.A(\mem[30] [2]), .B(\mem[31] [2]), .C(\adrram[0] ), 
         .Z(n1668)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1535_3_lut.init = 16'hcaca;
    LUT4 i1534_3_lut (.A(\mem[28] [2]), .B(\mem[29] [2]), .C(\adrram[0] ), 
         .Z(n1667)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1534_3_lut.init = 16'hcaca;
    LUT4 i1533_3_lut (.A(\mem[26] [2]), .B(\mem[27] [2]), .C(\adrram[0] ), 
         .Z(n1666)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1533_3_lut.init = 16'hcaca;
    LUT4 i1532_3_lut (.A(\mem[24] [2]), .B(\mem[25] [2]), .C(\adrram[0] ), 
         .Z(n1665)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1532_3_lut.init = 16'hcaca;
    LUT4 i1833_3_lut (.A(\mem[38] [3]), .B(\mem[39] [3]), .C(\adrram[0] ), 
         .Z(n1966)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1833_3_lut.init = 16'hcaca;
    LUT4 i1832_3_lut (.A(\mem[36] [3]), .B(\mem[37] [3]), .C(\adrram[0] ), 
         .Z(n1965)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1832_3_lut.init = 16'hcaca;
    LUT4 i1903_3_lut (.A(\mem[54] [1]), .B(\mem[55] [1]), .C(\adrram[0] ), 
         .Z(n2036)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1903_3_lut.init = 16'hcaca;
    LUT4 i1902_3_lut (.A(\mem[52] [1]), .B(\mem[53] [1]), .C(\adrram[0] ), 
         .Z(n2035)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1902_3_lut.init = 16'hcaca;
    LUT4 i1938_3_lut (.A(\mem[62] [0]), .B(\mem[63] [0]), .C(\adrram[0] ), 
         .Z(n2071)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1938_3_lut.init = 16'hcaca;
    LUT4 i1937_3_lut (.A(\mem[60] [0]), .B(\mem[61] [0]), .C(\adrram[0] ), 
         .Z(n2070)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1937_3_lut.init = 16'hcaca;
    LUT4 i1473_3_lut (.A(\mem[30] [0]), .B(\mem[31] [0]), .C(\adrram[0] ), 
         .Z(n1606)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1473_3_lut.init = 16'hcaca;
    LUT4 i1472_3_lut (.A(\mem[28] [0]), .B(\mem[29] [0]), .C(\adrram[0] ), 
         .Z(n1605)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1472_3_lut.init = 16'hcaca;
    LUT4 i1531_3_lut (.A(\mem[22] [2]), .B(\mem[23] [2]), .C(\adrram[0] ), 
         .Z(n1664)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1531_3_lut.init = 16'hcaca;
    LUT4 i1530_3_lut (.A(\mem[20] [2]), .B(\mem[21] [2]), .C(\adrram[0] ), 
         .Z(n1663)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1530_3_lut.init = 16'hcaca;
    LUT4 i1529_3_lut (.A(\mem[18] [2]), .B(\mem[19] [2]), .C(\adrram[0] ), 
         .Z(n1662)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1529_3_lut.init = 16'hcaca;
    LUT4 i1528_3_lut (.A(\mem[16] [2]), .B(\mem[17] [2]), .C(\adrram[0] ), 
         .Z(n1661)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1528_3_lut.init = 16'hcaca;
    LUT4 i1527_3_lut (.A(\mem[14] [2]), .B(\mem[15] [2]), .C(\adrram[0] ), 
         .Z(n1660)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1527_3_lut.init = 16'hcaca;
    LUT4 i1526_3_lut (.A(\mem[12] [2]), .B(\mem[13] [2]), .C(\adrram[0] ), 
         .Z(n1659)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1526_3_lut.init = 16'hcaca;
    LUT4 i1525_3_lut (.A(\mem[10] [2]), .B(\mem[11] [2]), .C(\adrram[0] ), 
         .Z(n1658)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1525_3_lut.init = 16'hcaca;
    LUT4 i1524_3_lut (.A(\mem[8] [2]), .B(\mem[9] [2]), .C(\adrram[0] ), 
         .Z(n1657)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1524_3_lut.init = 16'hcaca;
    LUT4 i1523_3_lut (.A(\mem[6] [2]), .B(\mem[7] [2]), .C(\adrram[0] ), 
         .Z(n1656)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1523_3_lut.init = 16'hcaca;
    LUT4 i1522_3_lut (.A(\mem[4] [2]), .B(\mem[5] [2]), .C(\adrram[0] ), 
         .Z(n1655)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1522_3_lut.init = 16'hcaca;
    LUT4 i1521_3_lut (.A(\mem[2] [2]), .B(\mem[3] [2]), .C(\adrram[0] ), 
         .Z(n1654)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1521_3_lut.init = 16'hcaca;
    LUT4 i1520_3_lut (.A(\mem[0] [2]), .B(\mem[1] [2]), .C(\adrram[0] ), 
         .Z(n1653)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1520_3_lut.init = 16'hcaca;
    LUT4 i2232_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2307), .C(n2306), 
         .D(\adrram[5] ), .Z(we_N_63_enable_224)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2232_2_lut_2_lut_3_lut_4_lut.init = 16'h0020;
    LUT4 i2287_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2307), .C(n2310), 
         .D(\adrram[5] ), .Z(we_N_63_enable_280)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2287_2_lut_2_lut_3_lut_4_lut.init = 16'h0002;
    LUT4 Select_672_i3_4_lut (.A(data_7__N_66[4]), .B(akku_o_c_4), .C(oe_N_57), 
         .D(n2305), .Z(data[4])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((D)+!B)) */ ;
    defparam Select_672_i3_4_lut.init = 16'ha0ec;
    LUT4 i2226_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2315), .C(n2306), 
         .D(\adrram[5] ), .Z(we_N_63_enable_216)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2226_2_lut_2_lut_3_lut_4_lut.init = 16'h0020;
    LUT4 i2299_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2315), .C(n2314), 
         .D(\adrram[5] ), .Z(we_N_63_enable_329)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2299_2_lut_2_lut_3_lut_4_lut.init = 16'h0002;
    LUT4 Select_673_i3_4_lut (.A(data_7__N_66[3]), .B(akku_o_c_3), .C(oe_N_57), 
         .D(n2305), .Z(data[3])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((D)+!B)) */ ;
    defparam Select_673_i3_4_lut.init = 16'ha0ec;
    LUT4 i2284_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2315), .C(n2310), 
         .D(\adrram[5] ), .Z(we_N_63_enable_273)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2284_2_lut_2_lut_3_lut_4_lut.init = 16'h0002;
    LUT4 i2246_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2309), .C(n2314), 
         .D(\adrram[5] ), .Z(we_N_63_enable_322)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2246_2_lut_2_lut_3_lut_4_lut.init = 16'h0002;
    LUT4 i2296_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2309), .C(n2306), 
         .D(\adrram[5] ), .Z(we_N_63_enable_201)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2296_2_lut_2_lut_3_lut_4_lut.init = 16'h0020;
    LUT4 i2281_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2309), .C(n2310), 
         .D(\adrram[5] ), .Z(we_N_63_enable_266)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2281_2_lut_2_lut_3_lut_4_lut.init = 16'h0002;
    LUT4 i1899_3_lut (.A(\mem[46] [1]), .B(\mem[47] [1]), .C(\adrram[0] ), 
         .Z(n2032)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1899_3_lut.init = 16'hcaca;
    LUT4 i2223_2_lut_2_lut_3_lut_4_lut (.A(\adrram[5] ), .B(n2308), .C(n2315), 
         .D(\adrram[2] ), .Z(we_N_63_enable_132)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2223_2_lut_2_lut_3_lut_4_lut.init = 16'h0200;
    LUT4 i2311_2_lut_2_lut_3_lut_4_lut (.A(\adrram[5] ), .B(n2308), .C(n2309), 
         .D(\adrram[2] ), .Z(we_N_63_enable_133)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2311_2_lut_2_lut_3_lut_4_lut.init = 16'h0200;
    LUT4 i2316_2_lut_2_lut_3_lut_4_lut (.A(\adrram[5] ), .B(n2308), .C(n2313), 
         .D(\adrram[2] ), .Z(we_N_63_enable_134)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2316_2_lut_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i2220_2_lut_2_lut_3_lut_4_lut (.A(\adrram[5] ), .B(n2308), .C(n2307), 
         .D(\adrram[2] ), .Z(we_N_63_enable_131)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2220_2_lut_2_lut_3_lut_4_lut.init = 16'h0200;
    LUT4 i2206_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2307), .C(n2314), 
         .D(\adrram[5] ), .Z(we_N_63_enable_368)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2206_2_lut_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i2345_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2307), .C(n2308), 
         .D(\adrram[5] ), .Z(we_N_63_enable_173)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2345_2_lut_2_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i2238_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2307), .C(n2310), 
         .D(\adrram[5] ), .Z(we_N_63_enable_308)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2238_2_lut_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i2276_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2307), .C(n2306), 
         .D(\adrram[5] ), .Z(we_N_63_enable_252)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2276_2_lut_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i2387_2_lut_2_lut_3_lut_4_lut (.A(\adrram[5] ), .B(n2308), .C(n2307), 
         .D(\adrram[2] ), .Z(we_N_63_enable_379)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2387_2_lut_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i2208_2_lut_2_lut_3_lut_4_lut (.A(\adrram[5] ), .B(n2308), .C(n2313), 
         .D(\adrram[2] ), .Z(we_N_63_enable_377)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2208_2_lut_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i2211_2_lut_2_lut_3_lut_4_lut (.A(\adrram[5] ), .B(n2308), .C(n2309), 
         .D(\adrram[2] ), .Z(we_N_63_enable_386)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2211_2_lut_2_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i2214_2_lut_2_lut_3_lut_4_lut (.A(\adrram[5] ), .B(n2308), .C(n2315), 
         .D(\adrram[2] ), .Z(we_N_63_enable_395)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2214_2_lut_2_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i2217_2_lut_2_lut_3_lut_4_lut (.A(\adrram[5] ), .B(n2308), .C(n2307), 
         .D(\adrram[2] ), .Z(we_N_63_enable_407)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2217_2_lut_2_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i1898_3_lut (.A(\mem[44] [1]), .B(\mem[45] [1]), .C(\adrram[0] ), 
         .Z(n2031)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1898_3_lut.init = 16'hcaca;
    LUT4 i2198_2_lut_2_lut_3_lut_4_lut (.A(\adrram[5] ), .B(n2310), .C(n2307), 
         .D(\adrram[2] ), .Z(we_N_63_enable_143)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2198_2_lut_2_lut_3_lut_4_lut.init = 16'h0002;
    LUT4 i2370_2_lut_2_lut_3_lut_4_lut (.A(\adrram[5] ), .B(n2310), .C(n2313), 
         .D(\adrram[2] ), .Z(we_N_63_enable_483)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2370_2_lut_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i2368_2_lut_2_lut_3_lut_4_lut (.A(\adrram[5] ), .B(n2310), .C(n2309), 
         .D(\adrram[2] ), .Z(we_N_63_enable_490)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2368_2_lut_2_lut_3_lut_4_lut.init = 16'h0200;
    LUT4 i2365_2_lut_2_lut_3_lut_4_lut (.A(\adrram[5] ), .B(n2310), .C(n2315), 
         .D(\adrram[2] ), .Z(we_N_63_enable_497)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2365_2_lut_2_lut_3_lut_4_lut.init = 16'h0200;
    LUT4 i2362_2_lut_2_lut_3_lut_4_lut (.A(\adrram[5] ), .B(n2310), .C(n2307), 
         .D(\adrram[2] ), .Z(we_N_63_enable_504)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2362_2_lut_2_lut_3_lut_4_lut.init = 16'h0200;
    LUT4 i2189_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2309), .C(n2314), 
         .D(\adrram[5] ), .Z(we_N_63_enable_351)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2189_2_lut_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i2340_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2309), .C(n2308), 
         .D(\adrram[5] ), .Z(we_N_63_enable_481)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2340_2_lut_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i2243_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2309), .C(n2306), 
         .D(\adrram[5] ), .Z(we_N_63_enable_238)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2243_2_lut_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i2195_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2309), .C(n2308), 
         .D(\adrram[5] ), .Z(we_N_63_enable_129)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2195_2_lut_2_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i2331_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2309), .C(n2310), 
         .D(\adrram[5] ), .Z(we_N_63_enable_512)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2331_2_lut_2_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i2293_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2309), .C(n2310), 
         .D(\adrram[5] ), .Z(we_N_63_enable_294)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2293_2_lut_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i2380_2_lut_2_lut_3_lut_4_lut (.A(\adrram[5] ), .B(n2306), .C(n2307), 
         .D(\adrram[2] ), .Z(we_N_63_enable_437)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i2380_2_lut_2_lut_3_lut_4_lut.init = 16'h0800;
    LUT4 i1164_2_lut_3_lut_4_lut (.A(\adrram[5] ), .B(n2306), .C(n2313), 
         .D(\adrram[2] ), .Z(we_N_63_enable_405)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1164_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i2376_2_lut_2_lut_3_lut_4_lut (.A(\adrram[5] ), .B(n2306), .C(n2309), 
         .D(\adrram[2] ), .Z(we_N_63_enable_455)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i2376_2_lut_2_lut_3_lut_4_lut.init = 16'h0008;
    LUT4 i2382_2_lut_2_lut_3_lut_4_lut (.A(\adrram[5] ), .B(n2306), .C(n2315), 
         .D(\adrram[2] ), .Z(we_N_63_enable_428)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i2382_2_lut_2_lut_3_lut_4_lut.init = 16'h0800;
    LUT4 i2384_2_lut_2_lut_3_lut_4_lut (.A(\adrram[5] ), .B(n2306), .C(n2309), 
         .D(\adrram[2] ), .Z(we_N_63_enable_420)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i2384_2_lut_2_lut_3_lut_4_lut.init = 16'h0800;
    LUT4 i2372_2_lut_2_lut_3_lut_4_lut (.A(\adrram[5] ), .B(n2306), .C(n2307), 
         .D(\adrram[2] ), .Z(we_N_63_enable_474)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i2372_2_lut_2_lut_3_lut_4_lut.init = 16'h0008;
    LUT4 i2328_2_lut_2_lut_3_lut_4_lut (.A(\adrram[5] ), .B(n2314), .C(n2309), 
         .D(\adrram[2] ), .Z(we_N_63_enable_137)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2328_2_lut_2_lut_3_lut_4_lut.init = 16'h0002;
    LUT4 i2319_2_lut_2_lut_3_lut_4_lut (.A(\adrram[5] ), .B(n2314), .C(n2307), 
         .D(\adrram[2] ), .Z(we_N_63_enable_135)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2319_2_lut_2_lut_3_lut_4_lut.init = 16'h0002;
    LUT4 i2356_2_lut_2_lut_3_lut_4_lut (.A(\adrram[5] ), .B(n2314), .C(n2313), 
         .D(\adrram[2] ), .Z(we_N_63_enable_174)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2356_2_lut_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i2354_2_lut_2_lut_3_lut_4_lut (.A(\adrram[5] ), .B(n2314), .C(n2309), 
         .D(\adrram[2] ), .Z(we_N_63_enable_188)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2354_2_lut_2_lut_3_lut_4_lut.init = 16'h0200;
    LUT4 i2351_2_lut_2_lut_3_lut_4_lut (.A(\adrram[5] ), .B(n2314), .C(n2315), 
         .D(\adrram[2] ), .Z(we_N_63_enable_202)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2351_2_lut_2_lut_3_lut_4_lut.init = 16'h0200;
    LUT4 i2348_2_lut_2_lut_3_lut_4_lut (.A(\adrram[5] ), .B(n2314), .C(n2307), 
         .D(\adrram[2] ), .Z(we_N_63_enable_213)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2348_2_lut_2_lut_3_lut_4_lut.init = 16'h0200;
    LUT4 i2325_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2313), .C(n2308), 
         .D(\adrram[5] ), .Z(we_N_63_enable_416)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2325_2_lut_2_lut_3_lut_4_lut.init = 16'h0004;
    LUT4 i669_1_lut (.A(\adrram[0] ), .Z(\pc_5__N_30[0] )) /* synthesis lut_function=(!(A)) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i669_1_lut.init = 16'h5555;
    LUT4 i1504_3_lut (.A(\mem[30] [1]), .B(\mem[31] [1]), .C(\adrram[0] ), 
         .Z(n1637)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1504_3_lut.init = 16'hcaca;
    LUT4 i1831_3_lut (.A(\mem[34] [3]), .B(\mem[35] [3]), .C(\adrram[0] ), 
         .Z(n1964)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1831_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_22 (.A(\adrram[0] ), .B(\adrram[1] ), .Z(n2309)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i1_2_lut_rep_22.init = 16'hbbbb;
    LUT4 i1_2_lut_rep_23 (.A(\adrram[3] ), .B(\adrram[4] ), .Z(n2310)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i1_2_lut_rep_23.init = 16'hbbbb;
    LUT4 i1_2_lut_rep_21 (.A(\adrram[3] ), .B(\adrram[4] ), .Z(n2308)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i1_2_lut_rep_21.init = 16'heeee;
    LUT4 i1830_3_lut (.A(\mem[32] [3]), .B(\mem[33] [3]), .C(\adrram[0] ), 
         .Z(n1963)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1830_3_lut.init = 16'hcaca;
    PFUMX i1912 (.BLUT(n2033), .ALUT(n2034), .C0(\adrram[1] ), .Z(n2045));
    L6MUX21 i1580 (.D0(n1710), .D1(n1711), .SD(\adrram[3] ), .Z(n1713));
    LUT4 i1_2_lut_rep_27 (.A(\adrram[4] ), .B(\adrram[3] ), .Z(n2314)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i1_2_lut_rep_27.init = 16'hbbbb;
    LUT4 i1503_3_lut (.A(\mem[28] [1]), .B(\mem[29] [1]), .C(\adrram[0] ), 
         .Z(n1636)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1503_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_28 (.A(\adrram[1] ), .B(\adrram[0] ), .Z(n2315)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i1_2_lut_rep_28.init = 16'hbbbb;
    L6MUX21 i1796 (.D0(n1925), .D1(n1926), .SD(\adrram[3] ), .Z(n1929));
    LUT4 i1936_3_lut (.A(\mem[58] [0]), .B(\mem[59] [0]), .C(\adrram[0] ), 
         .Z(n2069)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1936_3_lut.init = 16'hcaca;
    L6MUX21 i1797 (.D0(n1927), .D1(n1928), .SD(\adrram[3] ), .Z(n1930));
    L6MUX21 i1889 (.D0(n2018), .D1(n2019), .SD(\adrram[3] ), .Z(n2022));
    LUT4 i1935_3_lut (.A(\mem[56] [0]), .B(\mem[57] [0]), .C(\adrram[0] ), 
         .Z(n2068)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1935_3_lut.init = 16'hcaca;
    LUT4 Select_670_i3_4_lut (.A(data_7__N_66[6]), .B(akku_o_c_6), .C(oe_N_57), 
         .D(n2305), .Z(data[6])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((D)+!B)) */ ;
    defparam Select_670_i3_4_lut.init = 16'ha0ec;
    LUT4 i2235_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2313), .C(n2306), 
         .D(\adrram[5] ), .Z(we_N_63_enable_231)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2235_2_lut_2_lut_3_lut_4_lut.init = 16'h0040;
    L6MUX21 i1890 (.D0(n2020), .D1(n2021), .SD(\adrram[3] ), .Z(n2023));
    LUT4 i2201_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2313), .C(n2308), 
         .D(\adrram[5] ), .Z(we_N_63_enable_130)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2201_2_lut_2_lut_3_lut_4_lut.init = 16'h0400;
    LUT4 i2359_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2313), .C(n2310), 
         .D(\adrram[5] ), .Z(we_N_63_enable_511)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2359_2_lut_2_lut_3_lut_4_lut.init = 16'h0400;
    L6MUX21 i1641 (.D0(n1770), .D1(n1771), .SD(\adrram[3] ), .Z(n1774));
    LUT4 i1550_3_lut (.A(n1681), .B(n1682), .C(\adrram[4] ), .Z(n1683)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1550_3_lut.init = 16'hcaca;
    L6MUX21 i1642 (.D0(n1772), .D1(n1773), .SD(\adrram[3] ), .Z(n1775));
    LUT4 i1891_3_lut (.A(n2022), .B(n2023), .C(\adrram[4] ), .Z(n2024)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1891_3_lut.init = 16'hcaca;
    LUT4 Select_674_i3_4_lut (.A(data_7__N_66[2]), .B(akku_o_c_2), .C(oe_N_57), 
         .D(n2305), .Z(data[2])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((D)+!B)) */ ;
    defparam Select_674_i3_4_lut.init = 16'ha0ec;
    LUT4 i1860_3_lut (.A(n1991), .B(n1992), .C(\adrram[4] ), .Z(n1993)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1860_3_lut.init = 16'hcaca;
    LUT4 i1953_3_lut (.A(n2084), .B(n2085), .C(\adrram[4] ), .Z(n2086)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1953_3_lut.init = 16'hcaca;
    FD1P3AX mem_50__i0_i7 (.D(data[7]), .SP(we_N_63_enable_512), .CK(we_N_63), 
            .Q(\mem[50] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=47, LSE_RLINE=47 */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(56[9] 62[16])
    defparam mem_50__i0_i7.GSR = "ENABLED";
    LUT4 i1488_3_lut (.A(n1619), .B(n1620), .C(\adrram[4] ), .Z(n1621)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1488_3_lut.init = 16'hcaca;
    LUT4 i2305_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2313), .C(n2314), 
         .D(\adrram[5] ), .Z(we_N_63_enable_343)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2305_2_lut_2_lut_3_lut_4_lut.init = 16'h0004;
    L6MUX21 i1672 (.D0(n1801), .D1(n1802), .SD(\adrram[3] ), .Z(n1805));
    L6MUX21 i1673 (.D0(n1803), .D1(n1804), .SD(\adrram[3] ), .Z(n1806));
    LUT4 i1581_3_lut (.A(n1712), .B(n1713), .C(\adrram[4] ), .Z(n1714)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1581_3_lut.init = 16'hcaca;
    L6MUX21 i1827 (.D0(n1956), .D1(n1957), .SD(\adrram[3] ), .Z(n1960));
    L6MUX21 i1828 (.D0(n1958), .D1(n1959), .SD(\adrram[3] ), .Z(n1961));
    L6MUX21 i1703 (.D0(n1832), .D1(n1833), .SD(\adrram[3] ), .Z(n1836));
    L6MUX21 i1704 (.D0(n1834), .D1(n1835), .SD(\adrram[3] ), .Z(n1837));
    L6MUX21 i1544 (.D0(n1669), .D1(n1670), .SD(\adrram[2] ), .Z(n1677));
    L6MUX21 i1545 (.D0(n1671), .D1(n1672), .SD(\adrram[2] ), .Z(n1678));
    L6MUX21 i1546 (.D0(n1673), .D1(n1674), .SD(\adrram[2] ), .Z(n1679));
    L6MUX21 i1547 (.D0(n1675), .D1(n1676), .SD(\adrram[2] ), .Z(n1680));
    L6MUX21 i1484 (.D0(n1611), .D1(n1612), .SD(\adrram[2] ), .Z(n1617));
    L6MUX21 i1947 (.D0(n2072), .D1(n2073), .SD(\adrram[2] ), .Z(n2080));
    L6MUX21 i1485 (.D0(n1613), .D1(n1614), .SD(\adrram[2] ), .Z(n1618));
    L6MUX21 i1916 (.D0(n2041), .D1(n2042), .SD(\adrram[2] ), .Z(n2049));
    L6MUX21 i1854 (.D0(n1979), .D1(n1980), .SD(\adrram[2] ), .Z(n1987));
    L6MUX21 i1730 (.D0(n1855), .D1(n1856), .SD(\adrram[2] ), .Z(n1863));
    L6MUX21 i1948 (.D0(n2074), .D1(n2075), .SD(\adrram[2] ), .Z(n2081));
    L6MUX21 i1917 (.D0(n2043), .D1(n2044), .SD(\adrram[2] ), .Z(n2050));
    L6MUX21 i1855 (.D0(n1981), .D1(n1982), .SD(\adrram[2] ), .Z(n1988));
    L6MUX21 i1731 (.D0(n1857), .D1(n1858), .SD(\adrram[2] ), .Z(n1864));
    L6MUX21 i1732 (.D0(n1859), .D1(n1860), .SD(\adrram[2] ), .Z(n1865));
    L6MUX21 i1609 (.D0(n1737), .D1(n1738), .SD(\adrram[2] ), .Z(n1742));
    L6MUX21 i1608 (.D0(n1735), .D1(n1736), .SD(\adrram[2] ), .Z(n1741));
    L6MUX21 i1856 (.D0(n1983), .D1(n1984), .SD(\adrram[2] ), .Z(n1989));
    L6MUX21 i1733 (.D0(n1861), .D1(n1862), .SD(\adrram[2] ), .Z(n1866));
    L6MUX21 i1607 (.D0(n1733), .D1(n1734), .SD(\adrram[2] ), .Z(n1740));
    L6MUX21 i1606 (.D0(n1731), .D1(n1732), .SD(\adrram[2] ), .Z(n1739));
    L6MUX21 i1918 (.D0(n2045), .D1(n2046), .SD(\adrram[2] ), .Z(n2051));
    L6MUX21 i1857 (.D0(n1985), .D1(n1986), .SD(\adrram[2] ), .Z(n1990));
    L6MUX21 i1949 (.D0(n2076), .D1(n2077), .SD(\adrram[2] ), .Z(n2082));
    L6MUX21 i1919 (.D0(n2047), .D1(n2048), .SD(\adrram[2] ), .Z(n2052));
    L6MUX21 i1950 (.D0(n2078), .D1(n2079), .SD(\adrram[2] ), .Z(n2083));
    L6MUX21 i1513 (.D0(n1638), .D1(n1639), .SD(\adrram[2] ), .Z(n1646));
    L6MUX21 i1514 (.D0(n1640), .D1(n1641), .SD(\adrram[2] ), .Z(n1647));
    L6MUX21 i1515 (.D0(n1642), .D1(n1643), .SD(\adrram[2] ), .Z(n1648));
    L6MUX21 i1761 (.D0(n1886), .D1(n1887), .SD(\adrram[2] ), .Z(n1894));
    L6MUX21 i1762 (.D0(n1888), .D1(n1889), .SD(\adrram[2] ), .Z(n1895));
    L6MUX21 i1763 (.D0(n1890), .D1(n1891), .SD(\adrram[2] ), .Z(n1896));
    L6MUX21 i1764 (.D0(n1892), .D1(n1893), .SD(\adrram[2] ), .Z(n1897));
    L6MUX21 i1516 (.D0(n1644), .D1(n1645), .SD(\adrram[2] ), .Z(n1649));
    L6MUX21 i1575 (.D0(n1700), .D1(n1701), .SD(\adrram[2] ), .Z(n1708));
    L6MUX21 i1885 (.D0(n2010), .D1(n2011), .SD(\adrram[2] ), .Z(n2018));
    L6MUX21 i1576 (.D0(n1702), .D1(n1703), .SD(\adrram[2] ), .Z(n1709));
    L6MUX21 i1577 (.D0(n1704), .D1(n1705), .SD(\adrram[2] ), .Z(n1710));
    L6MUX21 i1792 (.D0(n1917), .D1(n1918), .SD(\adrram[2] ), .Z(n1925));
    L6MUX21 i1578 (.D0(n1706), .D1(n1707), .SD(\adrram[2] ), .Z(n1711));
    L6MUX21 i1886 (.D0(n2012), .D1(n2013), .SD(\adrram[2] ), .Z(n2019));
    L6MUX21 i1793 (.D0(n1919), .D1(n1920), .SD(\adrram[2] ), .Z(n1926));
    L6MUX21 i1794 (.D0(n1921), .D1(n1922), .SD(\adrram[2] ), .Z(n1927));
    L6MUX21 i1887 (.D0(n2014), .D1(n2015), .SD(\adrram[2] ), .Z(n2020));
    L6MUX21 i1795 (.D0(n1923), .D1(n1924), .SD(\adrram[2] ), .Z(n1928));
    L6MUX21 i1888 (.D0(n2016), .D1(n2017), .SD(\adrram[2] ), .Z(n2021));
    L6MUX21 i1637 (.D0(n1762), .D1(n1763), .SD(\adrram[2] ), .Z(n1770));
    L6MUX21 i1638 (.D0(n1764), .D1(n1765), .SD(\adrram[2] ), .Z(n1771));
    L6MUX21 i1639 (.D0(n1766), .D1(n1767), .SD(\adrram[2] ), .Z(n1772));
    L6MUX21 i1640 (.D0(n1768), .D1(n1769), .SD(\adrram[2] ), .Z(n1773));
    L6MUX21 i1823 (.D0(n1948), .D1(n1949), .SD(\adrram[2] ), .Z(n1956));
    L6MUX21 i1824 (.D0(n1950), .D1(n1951), .SD(\adrram[2] ), .Z(n1957));
    L6MUX21 i1825 (.D0(n1952), .D1(n1953), .SD(\adrram[2] ), .Z(n1958));
    L6MUX21 i1826 (.D0(n1954), .D1(n1955), .SD(\adrram[2] ), .Z(n1959));
    L6MUX21 i1668 (.D0(n1793), .D1(n1794), .SD(\adrram[2] ), .Z(n1801));
    L6MUX21 i1669 (.D0(n1795), .D1(n1796), .SD(\adrram[2] ), .Z(n1802));
    L6MUX21 i1670 (.D0(n1797), .D1(n1798), .SD(\adrram[2] ), .Z(n1803));
    L6MUX21 i1671 (.D0(n1799), .D1(n1800), .SD(\adrram[2] ), .Z(n1804));
    L6MUX21 i1483 (.D0(n1609), .D1(n1610), .SD(\adrram[2] ), .Z(n1616));
    L6MUX21 i1699 (.D0(n1824), .D1(n1825), .SD(\adrram[2] ), .Z(n1832));
    L6MUX21 i1700 (.D0(n1826), .D1(n1827), .SD(\adrram[2] ), .Z(n1833));
    L6MUX21 i1701 (.D0(n1828), .D1(n1829), .SD(\adrram[2] ), .Z(n1834));
    L6MUX21 i1702 (.D0(n1830), .D1(n1831), .SD(\adrram[2] ), .Z(n1835));
    L6MUX21 i1482 (.D0(n1607), .D1(n1608), .SD(\adrram[2] ), .Z(n1615));
    PFUMX i1536 (.BLUT(n1653), .ALUT(n1654), .C0(\adrram[1] ), .Z(n1669));
    PFUMX i1537 (.BLUT(n1655), .ALUT(n1656), .C0(\adrram[1] ), .Z(n1670));
    PFUMX i1538 (.BLUT(n1657), .ALUT(n1658), .C0(\adrram[1] ), .Z(n1671));
    PFUMX i1539 (.BLUT(n1659), .ALUT(n1660), .C0(\adrram[1] ), .Z(n1672));
    PFUMX i1540 (.BLUT(n1661), .ALUT(n1662), .C0(\adrram[1] ), .Z(n1673));
    PFUMX i1541 (.BLUT(n1663), .ALUT(n1664), .C0(\adrram[1] ), .Z(n1674));
    PFUMX i1481 (.BLUT(n1605), .ALUT(n1606), .C0(\adrram[1] ), .Z(n1614));
    PFUMX i1946 (.BLUT(n2070), .ALUT(n2071), .C0(\adrram[1] ), .Z(n2079));
    PFUMX i1913 (.BLUT(n2035), .ALUT(n2036), .C0(\adrram[1] ), .Z(n2046));
    PFUMX i1847 (.BLUT(n1965), .ALUT(n1966), .C0(\adrram[1] ), .Z(n1980));
    PFUMX i1542 (.BLUT(n1665), .ALUT(n1666), .C0(\adrram[1] ), .Z(n1675));
    PFUMX i1543 (.BLUT(n1667), .ALUT(n1668), .C0(\adrram[1] ), .Z(n1676));
    PFUMX i1848 (.BLUT(n1967), .ALUT(n1968), .C0(\adrram[1] ), .Z(n1981));
    PFUMX i1914 (.BLUT(n2037), .ALUT(n2038), .C0(\adrram[1] ), .Z(n2047));
    PFUMX i1849 (.BLUT(n1969), .ALUT(n1970), .C0(\adrram[1] ), .Z(n1982));
    PFUMX i1850 (.BLUT(n1971), .ALUT(n1972), .C0(\adrram[1] ), .Z(n1983));
    PFUMX i1722 (.BLUT(n1839), .ALUT(n1840), .C0(\adrram[1] ), .Z(n1855));
    PFUMX i1915 (.BLUT(n2039), .ALUT(n2040), .C0(\adrram[1] ), .Z(n2048));
    PFUMX i1851 (.BLUT(n1973), .ALUT(n1974), .C0(\adrram[1] ), .Z(n1984));
    PFUMX i1723 (.BLUT(n1841), .ALUT(n1842), .C0(\adrram[1] ), .Z(n1856));
    PFUMX i1724 (.BLUT(n1843), .ALUT(n1844), .C0(\adrram[1] ), .Z(n1857));
    PFUMX i1852 (.BLUT(n1975), .ALUT(n1976), .C0(\adrram[1] ), .Z(n1985));
    PFUMX i1725 (.BLUT(n1845), .ALUT(n1846), .C0(\adrram[1] ), .Z(n1858));
    PFUMX i1726 (.BLUT(n1847), .ALUT(n1848), .C0(\adrram[1] ), .Z(n1859));
    PFUMX i1754 (.BLUT(n1872), .ALUT(n1873), .C0(\adrram[1] ), .Z(n1887));
    PFUMX i1755 (.BLUT(n1874), .ALUT(n1875), .C0(\adrram[1] ), .Z(n1888));
    PFUMX i1756 (.BLUT(n1876), .ALUT(n1877), .C0(\adrram[1] ), .Z(n1889));
    PFUMX i1757 (.BLUT(n1878), .ALUT(n1879), .C0(\adrram[1] ), .Z(n1890));
    PFUMX i1758 (.BLUT(n1880), .ALUT(n1881), .C0(\adrram[1] ), .Z(n1891));
    PFUMX i1790 (.BLUT(n1913), .ALUT(n1914), .C0(\adrram[1] ), .Z(n1923));
    PFUMX i1505 (.BLUT(n1622), .ALUT(n1623), .C0(\adrram[1] ), .Z(n1638));
    PFUMX i1599 (.BLUT(n1717), .ALUT(n1718), .C0(\adrram[1] ), .Z(n1732));
    PFUMX i1506 (.BLUT(n1624), .ALUT(n1625), .C0(\adrram[1] ), .Z(n1639));
    PFUMX i1508 (.BLUT(n1628), .ALUT(n1629), .C0(\adrram[1] ), .Z(n1641));
    PFUMX i1883 (.BLUT(n2006), .ALUT(n2007), .C0(\adrram[1] ), .Z(n2016));
    PFUMX i1788 (.BLUT(n1909), .ALUT(n1910), .C0(\adrram[1] ), .Z(n1921));
    PFUMX i1509 (.BLUT(n1630), .ALUT(n1631), .C0(\adrram[1] ), .Z(n1642));
    PFUMX i1759 (.BLUT(n1882), .ALUT(n1883), .C0(\adrram[1] ), .Z(n1892));
    PFUMX i1760 (.BLUT(n1884), .ALUT(n1885), .C0(\adrram[1] ), .Z(n1893));
    PFUMX i1567 (.BLUT(n1684), .ALUT(n1685), .C0(\adrram[1] ), .Z(n1700));
    PFUMX i1568 (.BLUT(n1686), .ALUT(n1687), .C0(\adrram[1] ), .Z(n1701));
    PFUMX i1884 (.BLUT(n2008), .ALUT(n2009), .C0(\adrram[1] ), .Z(n2017));
    PFUMX i1789 (.BLUT(n1911), .ALUT(n1912), .C0(\adrram[1] ), .Z(n1922));
    PFUMX i1753 (.BLUT(n1870), .ALUT(n1871), .C0(\adrram[1] ), .Z(n1886));
    PFUMX i1474 (.BLUT(n1591), .ALUT(n1592), .C0(\adrram[1] ), .Z(n1607));
    PFUMX i1600 (.BLUT(n1719), .ALUT(n1720), .C0(\adrram[1] ), .Z(n1733));
    PFUMX i1601 (.BLUT(n1721), .ALUT(n1722), .C0(\adrram[1] ), .Z(n1734));
    PFUMX i1602 (.BLUT(n1723), .ALUT(n1724), .C0(\adrram[1] ), .Z(n1735));
    PFUMX i1603 (.BLUT(n1725), .ALUT(n1726), .C0(\adrram[1] ), .Z(n1736));
    PFUMX i1604 (.BLUT(n1727), .ALUT(n1728), .C0(\adrram[1] ), .Z(n1737));
    PFUMX i1605 (.BLUT(n1729), .ALUT(n1730), .C0(\adrram[1] ), .Z(n1738));
    PFUMX i1729 (.BLUT(n1853), .ALUT(n1854), .C0(\adrram[1] ), .Z(n1862));
    PFUMX i1728 (.BLUT(n1851), .ALUT(n1852), .C0(\adrram[1] ), .Z(n1861));
    PFUMX i1727 (.BLUT(n1849), .ALUT(n1850), .C0(\adrram[1] ), .Z(n1860));
    PFUMX i1853 (.BLUT(n1977), .ALUT(n1978), .C0(\adrram[1] ), .Z(n1986));
    PFUMX i1569 (.BLUT(n1688), .ALUT(n1689), .C0(\adrram[1] ), .Z(n1702));
    PFUMX i1787 (.BLUT(n1907), .ALUT(n1908), .C0(\adrram[1] ), .Z(n1920));
    PFUMX i1660 (.BLUT(n1777), .ALUT(n1778), .C0(\adrram[1] ), .Z(n1793));
    PFUMX i1480 (.BLUT(n1603), .ALUT(n1604), .C0(\adrram[1] ), .Z(n1613));
    PFUMX i1629 (.BLUT(n1746), .ALUT(n1747), .C0(\adrram[1] ), .Z(n1762));
    PFUMX i1634 (.BLUT(n1756), .ALUT(n1757), .C0(\adrram[1] ), .Z(n1767));
    PFUMX i1939 (.BLUT(n2056), .ALUT(n2057), .C0(\adrram[1] ), .Z(n2072));
    PFUMX i1691 (.BLUT(n1808), .ALUT(n1809), .C0(\adrram[1] ), .Z(n1824));
    PFUMX i1661 (.BLUT(n1779), .ALUT(n1780), .C0(\adrram[1] ), .Z(n1794));
    PFUMX i1510 (.BLUT(n1632), .ALUT(n1633), .C0(\adrram[1] ), .Z(n1643));
    PFUMX i1692 (.BLUT(n1810), .ALUT(n1811), .C0(\adrram[1] ), .Z(n1825));
    PFUMX i1662 (.BLUT(n1781), .ALUT(n1782), .C0(\adrram[1] ), .Z(n1795));
    PFUMX i1630 (.BLUT(n1748), .ALUT(n1749), .C0(\adrram[1] ), .Z(n1763));
    PFUMX i1635 (.BLUT(n1758), .ALUT(n1759), .C0(\adrram[1] ), .Z(n1768));
    PFUMX i1818 (.BLUT(n1938), .ALUT(n1939), .C0(\adrram[1] ), .Z(n1951));
    PFUMX i1693 (.BLUT(n1812), .ALUT(n1813), .C0(\adrram[1] ), .Z(n1826));
    PFUMX i1663 (.BLUT(n1783), .ALUT(n1784), .C0(\adrram[1] ), .Z(n1796));
    PFUMX i1791 (.BLUT(n1915), .ALUT(n1916), .C0(\adrram[1] ), .Z(n1924));
    PFUMX i1694 (.BLUT(n1814), .ALUT(n1815), .C0(\adrram[1] ), .Z(n1827));
    PFUMX i1664 (.BLUT(n1785), .ALUT(n1786), .C0(\adrram[1] ), .Z(n1797));
    PFUMX i1636 (.BLUT(n1760), .ALUT(n1761), .C0(\adrram[1] ), .Z(n1769));
    PFUMX i1819 (.BLUT(n1940), .ALUT(n1941), .C0(\adrram[1] ), .Z(n1952));
    PFUMX i1695 (.BLUT(n1816), .ALUT(n1817), .C0(\adrram[1] ), .Z(n1828));
    PFUMX i1665 (.BLUT(n1787), .ALUT(n1788), .C0(\adrram[1] ), .Z(n1798));
    PFUMX i1696 (.BLUT(n1818), .ALUT(n1819), .C0(\adrram[1] ), .Z(n1829));
    PFUMX i1666 (.BLUT(n1789), .ALUT(n1790), .C0(\adrram[1] ), .Z(n1799));
    PFUMX i1820 (.BLUT(n1942), .ALUT(n1943), .C0(\adrram[1] ), .Z(n1953));
    PFUMX i1909 (.BLUT(n2027), .ALUT(n2028), .C0(\adrram[1] ), .Z(n2042));
    PFUMX i1941 (.BLUT(n2060), .ALUT(n2061), .C0(\adrram[1] ), .Z(n2074));
    PFUMX i1631 (.BLUT(n1750), .ALUT(n1751), .C0(\adrram[1] ), .Z(n1764));
    LUT4 i1829_3_lut (.A(n1960), .B(n1961), .C(\adrram[4] ), .Z(n1962)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1829_3_lut.init = 16'hcaca;
    PFUMX i1511 (.BLUT(n1634), .ALUT(n1635), .C0(\adrram[1] ), .Z(n1644));
    PFUMX i1815 (.BLUT(n1932), .ALUT(n1933), .C0(\adrram[1] ), .Z(n1948));
    PFUMX i1910 (.BLUT(n2029), .ALUT(n2030), .C0(\adrram[1] ), .Z(n2043));
    LUT4 i2334_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2313), .C(n2314), 
         .D(\adrram[5] ), .Z(we_N_63_enable_219)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2334_2_lut_2_lut_3_lut_4_lut.init = 16'h0400;
    PFUMX i1507 (.BLUT(n1626), .ALUT(n1627), .C0(\adrram[1] ), .Z(n1640));
    PFUMX i1598 (.BLUT(n1715), .ALUT(n1716), .C0(\adrram[1] ), .Z(n1731));
    PFUMX i1821 (.BLUT(n1944), .ALUT(n1945), .C0(\adrram[1] ), .Z(n1954));
    PFUMX i1667 (.BLUT(n1791), .ALUT(n1792), .C0(\adrram[1] ), .Z(n1800));
    LUT4 i1612_3_lut (.A(n1743), .B(n1744), .C(\adrram[4] ), .Z(n1745)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1612_3_lut.init = 16'hcaca;
    PFUMX i1632 (.BLUT(n1752), .ALUT(n1753), .C0(\adrram[1] ), .Z(n1765));
    PFUMX i1816 (.BLUT(n1934), .ALUT(n1935), .C0(\adrram[1] ), .Z(n1949));
    PFUMX i1697 (.BLUT(n1820), .ALUT(n1821), .C0(\adrram[1] ), .Z(n1830));
    LUT4 Select_675_i3_4_lut (.A(data_7__N_66[1]), .B(akku_o_c_1), .C(oe_N_57), 
         .D(n2305), .Z(data[1])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((D)+!B)) */ ;
    defparam Select_675_i3_4_lut.init = 16'ha0ec;
    PFUMX i1940 (.BLUT(n2058), .ALUT(n2059), .C0(\adrram[1] ), .Z(n2073));
    PFUMX i1942 (.BLUT(n2062), .ALUT(n2063), .C0(\adrram[1] ), .Z(n2075));
    LUT4 i2290_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2313), .C(n2310), 
         .D(\adrram[5] ), .Z(we_N_63_enable_287)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2290_2_lut_2_lut_3_lut_4_lut.init = 16'h0004;
    LUT4 i1798_3_lut (.A(n1929), .B(n1930), .C(\adrram[4] ), .Z(n1931)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1798_3_lut.init = 16'hcaca;
    PFUMX i1633 (.BLUT(n1754), .ALUT(n1755), .C0(\adrram[1] ), .Z(n1766));
    PFUMX i1817 (.BLUT(n1936), .ALUT(n1937), .C0(\adrram[1] ), .Z(n1950));
    PFUMX i1944 (.BLUT(n2066), .ALUT(n2067), .C0(\adrram[1] ), .Z(n2077));
    LUT4 i1643_3_lut (.A(n1774), .B(n1775), .C(\adrram[4] ), .Z(n1776)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1643_3_lut.init = 16'hcaca;
    PFUMX i1822 (.BLUT(n1946), .ALUT(n1947), .C0(\adrram[1] ), .Z(n1955));
    PFUMX i1943 (.BLUT(n2064), .ALUT(n2065), .C0(\adrram[1] ), .Z(n2076));
    LUT4 i1767_3_lut (.A(n1898), .B(n1899), .C(\adrram[4] ), .Z(n1900)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1767_3_lut.init = 16'hcaca;
    LUT4 i1674_3_lut (.A(n1805), .B(n1806), .C(\adrram[4] ), .Z(n1807)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1674_3_lut.init = 16'hcaca;
    PFUMX i1698 (.BLUT(n1822), .ALUT(n1823), .C0(\adrram[1] ), .Z(n1831));
    LUT4 i1736_3_lut (.A(n1867), .B(n1868), .C(\adrram[4] ), .Z(n1869)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1736_3_lut.init = 16'hcaca;
    PFUMX i1908 (.BLUT(n2025), .ALUT(n2026), .C0(\adrram[1] ), .Z(n2041));
    PFUMX i1570 (.BLUT(n1690), .ALUT(n1691), .C0(\adrram[1] ), .Z(n1703));
    PFUMX i1571 (.BLUT(n1692), .ALUT(n1693), .C0(\adrram[1] ), .Z(n1704));
    PFUMX i1572 (.BLUT(n1694), .ALUT(n1695), .C0(\adrram[1] ), .Z(n1705));
    PFUMX i1573 (.BLUT(n1696), .ALUT(n1697), .C0(\adrram[1] ), .Z(n1706));
    PFUMX i1475 (.BLUT(n1593), .ALUT(n1594), .C0(\adrram[1] ), .Z(n1608));
    PFUMX i1574 (.BLUT(n1698), .ALUT(n1699), .C0(\adrram[1] ), .Z(n1707));
    PFUMX i1476 (.BLUT(n1595), .ALUT(n1596), .C0(\adrram[1] ), .Z(n1609));
    PFUMX i1477 (.BLUT(n1597), .ALUT(n1598), .C0(\adrram[1] ), .Z(n1610));
    PFUMX i1478 (.BLUT(n1599), .ALUT(n1600), .C0(\adrram[1] ), .Z(n1611));
    PFUMX i1877 (.BLUT(n1994), .ALUT(n1995), .C0(\adrram[1] ), .Z(n2010));
    PFUMX i1878 (.BLUT(n1996), .ALUT(n1997), .C0(\adrram[1] ), .Z(n2011));
    PFUMX i1479 (.BLUT(n1601), .ALUT(n1602), .C0(\adrram[1] ), .Z(n1612));
    PFUMX i1879 (.BLUT(n1998), .ALUT(n1999), .C0(\adrram[1] ), .Z(n2012));
    PFUMX i1880 (.BLUT(n2000), .ALUT(n2001), .C0(\adrram[1] ), .Z(n2013));
    PFUMX i1881 (.BLUT(n2002), .ALUT(n2003), .C0(\adrram[1] ), .Z(n2014));
    PFUMX i1784 (.BLUT(n1901), .ALUT(n1902), .C0(\adrram[1] ), .Z(n1917));
    PFUMX i1882 (.BLUT(n2004), .ALUT(n2005), .C0(\adrram[1] ), .Z(n2015));
    PFUMX i1785 (.BLUT(n1903), .ALUT(n1904), .C0(\adrram[1] ), .Z(n1918));
    LUT4 i1705_3_lut (.A(n1836), .B(n1837), .C(\adrram[4] ), .Z(n1838)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1705_3_lut.init = 16'hcaca;
    LUT4 Select_669_i3_4_lut (.A(data_7__N_66[7]), .B(akku_o_c_7), .C(oe_N_57), 
         .D(n2305), .Z(data[7])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((D)+!B)) */ ;
    defparam Select_669_i3_4_lut.init = 16'ha0ec;
    LUT4 i2378_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2313), .C(n2306), 
         .D(\adrram[5] ), .Z(we_N_63_enable_446)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2378_2_lut_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 i1901_3_lut (.A(\mem[50] [1]), .B(\mem[51] [1]), .C(\adrram[0] ), 
         .Z(n2034)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1901_3_lut.init = 16'hcaca;
    LUT4 i1690_3_lut (.A(\mem[30] [7]), .B(\mem[31] [7]), .C(\adrram[0] ), 
         .Z(n1823)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1690_3_lut.init = 16'hcaca;
    LUT4 i2337_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2315), .C(n2308), 
         .D(\adrram[5] ), .Z(we_N_63_enable_452)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2337_2_lut_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i2273_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2315), .C(n2306), 
         .D(\adrram[5] ), .Z(we_N_63_enable_245)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2273_2_lut_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i2308_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2315), .C(n2314), 
         .D(\adrram[5] ), .Z(we_N_63_enable_359)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2308_2_lut_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i2322_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2315), .C(n2314), 
         .D(\adrram[5] ), .Z(we_N_63_enable_136)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2322_2_lut_2_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i2192_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2315), .C(n2308), 
         .D(\adrram[5] ), .Z(we_N_63_enable_160)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2192_2_lut_2_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i2374_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2315), .C(n2306), 
         .D(\adrram[5] ), .Z(we_N_63_enable_465)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2374_2_lut_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i2229_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2315), .C(n2310), 
         .D(\adrram[5] ), .Z(we_N_63_enable_301)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2229_2_lut_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i2314_2_lut_2_lut_3_lut_4_lut (.A(\adrram[2] ), .B(n2315), .C(n2310), 
         .D(\adrram[5] ), .Z(we_N_63_enable_144)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i2314_2_lut_2_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i1155_2_lut_rep_19 (.A(\adrram[4] ), .B(\adrram[3] ), .Z(n2306)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1155_2_lut_rep_19.init = 16'h8888;
    LUT4 i1900_3_lut (.A(\mem[48] [1]), .B(\mem[49] [1]), .C(\adrram[0] ), 
         .Z(n2033)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1900_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_20 (.A(\adrram[1] ), .B(\adrram[0] ), .Z(n2307)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/70735/desktop/cpu/sram64kx8.vhd(60[21:47])
    defparam i1_2_lut_rep_20.init = 16'heeee;
    LUT4 i1922_3_lut (.A(n2053), .B(n2054), .C(\adrram[4] ), .Z(n2055)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1922_3_lut.init = 16'hcaca;
    LUT4 i1519_3_lut (.A(n1650), .B(n1651), .C(\adrram[4] ), .Z(n1652)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1519_3_lut.init = 16'hcaca;
    PFUMX i1786 (.BLUT(n1905), .ALUT(n1906), .C0(\adrram[1] ), .Z(n1919));
    
endmodule
//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

